VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 2000 ;
END UNITS

PROPERTYDEFINITIONS
    LAYER LEF58_CORNERSPACING STRING ;
END PROPERTYDEFINITIONS

CLEARANCEMEASURE EUCLIDEAN ;
MANUFACTURINGGRID 0.0005 ;
USEMINSPACING OBS ON ;

LAYER Metal1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.10 0.10 ;
  WIDTH 0.05 ;
  MINWIDTH 0.05 ;
  AREA 0.0115 ;
  SPACINGTABLE
    PARALLELRUNLENGTH  0.0 0.22 0.47 0.63 1.50
    WIDTH 0.0         0.05 0.05 0.05 0.05 0.05
    WIDTH 0.10        0.05 0.06 0.06 0.06 0.06
    WIDTH 0.28        0.05 0.10 0.10 0.10 0.10
    WIDTH 0.47        0.05 0.10 0.13 0.13 0.13
    WIDTH 0.63        0.05 0.10 0.13 0.15 0.15
    WIDTH 1.50        0.05 0.10 0.13 0.15 0.50 ;
  SPACING 0.06 ENDOFLINE 0.06 WITHIN 0.025 ;
END Metal1

LAYER Via1
  TYPE CUT ;
  SPACING 0.075 ;
  WIDTH 0.05 ;
END Via1

LAYER Metal2
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.10 0.10 ;
  WIDTH 0.05 ;
  MINWIDTH 0.05 ;
  AREA 0.014 ;
  SPACINGTABLE
    PARALLELRUNLENGTH  0.0 0.22 0.47 0.63 1.5
    WIDTH 0.0         0.05 0.05 0.05 0.05 0.05
    WIDTH 0.09        0.05 0.06 0.06 0.06 0.06
    WIDTH 0.16        0.05 0.10 0.10 0.10 0.10
    WIDTH 0.47        0.05 0.10 0.13 0.13 0.13
    WIDTH 0.63        0.05 0.10 0.13 0.15 0.15
    WIDTH 1.5         0.05 0.10 0.13 0.15 0.50 ;
  SPACING 0.08 ENDOFLINE 0.08 WITHIN 0.025 ;
  SPACING 0.10 ENDOFLINE 0.08 WITHIN 0.025 PARALLELEDGE 0.10 WITHIN 0.025 ;
  PROPERTY LEF58_CORNERSPACING "CORNERSPACING CONVEXCORNER EXCEPTEOL 0.08
    WIDTH 0.00 SPACING 0.10
    WIDTH 0.20 SPACING 0.20
    WIDTH 0.50 SPACING 0.30 ;" ;
END Metal2

LAYER Via2
  TYPE CUT ;
  SPACING 0.075 ;
  WIDTH 0.05 ;
  SPACING 0.155 ADJACENTCUTS 3 WITHIN 0.200 ;
END Via2

LAYER Metal3
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.10 0.10 ;
  WIDTH 0.05 ;
  MINWIDTH 0.05 ;
  AREA 0.017 ;
  SPACINGTABLE
    PARALLELRUNLENGTH  0.0 0.22 0.47 0.63 1.5
    WIDTH 0.0         0.05 0.05 0.05 0.05 0.05
    WIDTH 0.09        0.05 0.06 0.06 0.06 0.06
    WIDTH 0.16        0.05 0.10 0.10 0.10 0.10
    WIDTH 0.47        0.05 0.10 0.13 0.13 0.13
    WIDTH 0.63        0.05 0.10 0.13 0.15 0.15
    WIDTH 1.5         0.05 0.10 0.13 0.15 0.50 ;
  SPACING 0.08 ENDOFLINE 0.08 WITHIN 0.025 ;
  SPACING 0.10 ENDOFLINE 0.08 WITHIN 0.025 PARALLELEDGE 0.10 WITHIN 0.025 ;
  PROPERTY LEF58_CORNERSPACING "CORNERSPACING CONVEXCORNER EXCEPTEOL 0.08
    WIDTH 0.00 SPACING 0.10
    WIDTH 0.20 SPACING 0.20
    WIDTH 0.50 SPACING 0.30 ;" ;
END Metal3

LAYER Via3
  TYPE CUT ;
  SPACING 0.075 ;
  WIDTH 0.05 ;
  SPACING 0.155 ADJACENTCUTS 3 WITHIN 0.200 ;
END Via3

LAYER Metal4
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.10 0.10 ;
  WIDTH 0.05 ;
  MINWIDTH 0.05 ;
  AREA 0.017 ;
  SPACINGTABLE
    PARALLELRUNLENGTH  0.0 0.22 0.47 0.63 1.5
    WIDTH 0.0         0.05 0.05 0.05 0.05 0.05
    WIDTH 0.09        0.05 0.06 0.06 0.06 0.06
    WIDTH 0.16        0.05 0.10 0.10 0.10 0.10
    WIDTH 0.47        0.05 0.10 0.13 0.13 0.13
    WIDTH 0.63        0.05 0.10 0.13 0.15 0.15
    WIDTH 1.5         0.05 0.10 0.13 0.15 0.50 ;
  SPACING 0.08 ENDOFLINE 0.08 WITHIN 0.025 ;
  SPACING 0.10 ENDOFLINE 0.08 WITHIN 0.025 PARALLELEDGE 0.10 WITHIN 0.025 ;
  PROPERTY LEF58_CORNERSPACING "CORNERSPACING CONVEXCORNER EXCEPTEOL 0.08
    WIDTH 0.00 SPACING 0.10
    WIDTH 0.20 SPACING 0.20
    WIDTH 0.50 SPACING 0.30 ;" ;
END Metal4

LAYER Via4
  TYPE CUT ;
  SPACING 0.075 ;
  WIDTH 0.05 ;
  SPACING 0.155 ADJACENTCUTS 3 WITHIN 0.200 ;
END Via4

LAYER Metal5
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.10 0.10 ;
  WIDTH 0.05 ;
  MINWIDTH 0.05 ;
  AREA 0.017 ;
  SPACINGTABLE
    PARALLELRUNLENGTH  0.0 0.22 0.47 0.63 1.5
    WIDTH 0.0         0.05 0.05 0.05 0.05 0.05
    WIDTH 0.09        0.05 0.06 0.06 0.06 0.06
    WIDTH 0.16        0.05 0.10 0.10 0.10 0.10
    WIDTH 0.47        0.05 0.10 0.13 0.13 0.13
    WIDTH 0.63        0.05 0.10 0.13 0.15 0.15
    WIDTH 1.5         0.05 0.10 0.13 0.15 0.50 ;
  SPACING 0.08 ENDOFLINE 0.08 WITHIN 0.025 ;
  SPACING 0.10 ENDOFLINE 0.08 WITHIN 0.025 PARALLELEDGE 0.10 WITHIN 0.025 ;
  PROPERTY LEF58_CORNERSPACING "CORNERSPACING CONVEXCORNER EXCEPTEOL 0.08
    WIDTH 0.00 SPACING 0.10
    WIDTH 0.20 SPACING 0.20
    WIDTH 0.50 SPACING 0.30 ;" ;
END Metal5

LAYER Via5
  TYPE CUT ;
  SPACING 0.075 ;
  WIDTH 0.05 ;
  SPACING 0.155 ADJACENTCUTS 3 WITHIN 0.200 ;
END Via5

LAYER Metal6
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.15 0.15 ;
  WIDTH 0.07 ;
  MINWIDTH 0.07 ;
  AREA 0.025 ;
  SPACINGTABLE
    PARALLELRUNLENGTH  0.0 0.22 0.47 0.63 1.5
    WIDTH 0.0         0.08 0.08 0.08 0.08 0.08
    WIDTH 0.10        0.08 0.12 0.12 0.12 0.12
    WIDTH 0.16        0.08 0.12 0.15 0.15 0.15
    WIDTH 0.47        0.08 0.12 0.15 0.18 0.18
    WIDTH 0.63        0.08 0.12 0.15 0.18 0.25
    WIDTH 1.5         0.08 0.12 0.15 0.18 0.50 ;
  SPACING 0.10 ENDOFLINE 0.10 WITHIN 0.035 ;
  SPACING 0.12 ENDOFLINE 0.10 WITHIN 0.035 PARALLELEDGE 0.12 WITHIN 0.035 ;
  PROPERTY LEF58_CORNERSPACING "CORNERSPACING CONVEXCORNER EXCEPTEOL 0.08
    WIDTH 0.00 SPACING 0.10
    WIDTH 0.20 SPACING 0.20
    WIDTH 0.50 SPACING 0.30 ;" ;
END Metal6

LAYER Via6
  TYPE CUT ;
  SPACING 0.10 ;
  WIDTH 0.07 ;
  SPACING 0.20 ADJACENTCUTS 3 WITHIN 0.25 ;
END Via6

LAYER Metal7
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.15 0.15 ;
  WIDTH 0.07 ;
  MINWIDTH 0.07 ;
  AREA 0.025 ;
  SPACINGTABLE
    PARALLELRUNLENGTH  0.0 0.22 0.47 0.63 1.5
    WIDTH 0.0         0.08 0.08 0.08 0.08 0.08
    WIDTH 0.10        0.08 0.12 0.12 0.12 0.12
    WIDTH 0.16        0.08 0.12 0.15 0.15 0.15
    WIDTH 0.47        0.08 0.12 0.15 0.18 0.18
    WIDTH 0.63        0.08 0.12 0.15 0.18 0.25
    WIDTH 1.5         0.08 0.12 0.15 0.18 0.50 ;
  SPACING 0.10 ENDOFLINE 0.10 WITHIN 0.035 ;
  SPACING 0.12 ENDOFLINE 0.10 WITHIN 0.035 PARALLELEDGE 0.12 WITHIN 0.035 ;
  PROPERTY LEF58_CORNERSPACING "CORNERSPACING CONVEXCORNER EXCEPTEOL 0.08
    WIDTH 0.00 SPACING 0.10
    WIDTH 0.20 SPACING 0.20
    WIDTH 0.50 SPACING 0.30 ;" ;
END Metal7

LAYER Via7
  TYPE CUT ;
  SPACING 0.10 ;
  WIDTH 0.07 ;
  SPACING 0.20 ADJACENTCUTS 3 WITHIN 0.25 ;
END Via7

LAYER Metal8
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.2 0.2 ;
  WIDTH 0.10 ;
  MINWIDTH 0.10 ;
  AREA 0.052 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0.0 0.22 0.47 0.63 1.5
    WIDTH 0	     0.10 0.10 0.10 0.10 0.10
    WIDTH 0.2	     0.10 0.15 0.15 0.15 0.15
    WIDTH 0.4	     0.10 0.15 0.20 0.20 0.20
    WIDTH 1.5	     0.10 0.15 0.20 0.30 0.50 ;
  SPACING 0.12 ENDOFLINE 0.12 WITHIN 0.035 ;
END Metal8

LAYER Via8
  TYPE CUT ;
  SPACING 0.15 ;
  WIDTH 0.10 ;
END Via8

LAYER Metal9
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.2 0.2 ;
  WIDTH 0.10 ;
  MINWIDTH 0.10 ;
  AREA 0.052 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0.0 0.22 0.47 0.63 1.5
    WIDTH 0	     0.10 0.10 0.10 0.10 0.10
    WIDTH 0.2	     0.10 0.15 0.15 0.15 0.15
    WIDTH 0.4	     0.10 0.15 0.20 0.20 0.20
    WIDTH 1.5	     0.10 0.15 0.20 0.30 0.50 ;
  SPACING 0.12 ENDOFLINE 0.12 WITHIN 0.035 ;
END Metal9

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA VIA12_1C DEFAULT 
    LAYER Metal1 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
    LAYER Via1 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal2 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
END VIA12_1C

VIA VIA12_1C_H DEFAULT 
    LAYER Metal1 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
    LAYER Via1 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal2 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
END VIA12_1C_H

VIA VIA12_1C_V DEFAULT 
    LAYER Metal1 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
    LAYER Via1 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal2 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
END VIA12_1C_V

VIA VIA12_PG
    LAYER Metal1 ;
        RECT -0.350000 -0.050000 0.350000 0.050000 ;
    LAYER Via1 ;
        RECT -0.325000 -0.025000 -0.275000 0.025000 ;
        RECT -0.175000 -0.025000 -0.125000 0.025000 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
        RECT 0.125000 -0.025000 0.175000 0.025000 ;
        RECT 0.275000 -0.025000 0.325000 0.025000 ;
    LAYER Metal2 ;
        RECT -0.350000 -0.050000 0.350000 0.050000 ;
END VIA12_PG

VIA VIA23_1C DEFAULT 
    LAYER Metal2 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
    LAYER Via2 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal3 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
END VIA23_1C

VIA VIA23_1C_H DEFAULT 
    LAYER Metal2 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
    LAYER Via2 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal3 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
END VIA23_1C_H

VIA VIA23_1C_V DEFAULT 
    LAYER Metal2 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
    LAYER Via2 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal3 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
END VIA23_1C_V

VIA VIA23_1ST_E DEFAULT 
    LAYER Metal2 ;
        RECT -0.055000 -0.025000 0.325000 0.025000 ;
    LAYER Via2 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal3 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
END VIA23_1ST_E

VIA VIA23_1ST_W DEFAULT 
    LAYER Metal2 ;
        RECT -0.325000 -0.025000 0.055000 0.025000 ;
    LAYER Via2 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal3 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
END VIA23_1ST_W

VIA VIA23_PG
    LAYER Metal2 ;
        RECT -0.350000 -0.050000 0.350000 0.050000 ;
    LAYER Via2 ;
        RECT -0.325000 -0.025000 -0.275000 0.025000 ;
        RECT -0.175000 -0.025000 -0.125000 0.025000 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
        RECT 0.125000 -0.025000 0.175000 0.025000 ;
        RECT 0.275000 -0.025000 0.325000 0.025000 ;
    LAYER Metal3 ;
        RECT -0.350000 -0.050000 0.350000 0.050000 ;
END VIA23_PG

VIA VIA34_1C DEFAULT 
    LAYER Metal3 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
    LAYER Via3 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal4 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
END VIA34_1C

VIA VIA34_1C_H DEFAULT 
    LAYER Metal3 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
    LAYER Via3 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal4 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
END VIA34_1C_H

VIA VIA34_1C_V DEFAULT 
    LAYER Metal3 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
    LAYER Via3 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal4 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
END VIA34_1C_V

VIA VIA34_1ST_N DEFAULT 
    LAYER Metal3 ;
        RECT -0.025000 -0.055000 0.025000 0.325000 ;
    LAYER Via3 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal4 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
END VIA34_1ST_N

VIA VIA34_1ST_S DEFAULT 
    LAYER Metal3 ;
        RECT -0.025000 -0.325000 0.025000 0.055000 ;
    LAYER Via3 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal4 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
END VIA34_1ST_S

VIA VIA34_PG
    LAYER Metal3 ;
        RECT -0.350000 -0.050000 0.350000 0.050000 ;
    LAYER Via3 ;
        RECT -0.325000 -0.025000 -0.275000 0.025000 ;
        RECT -0.175000 -0.025000 -0.125000 0.025000 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
        RECT 0.125000 -0.025000 0.175000 0.025000 ;
        RECT 0.275000 -0.025000 0.325000 0.025000 ;
    LAYER Metal4 ;
        RECT -0.350000 -0.050000 0.350000 0.050000 ;
END VIA34_PG

VIA VIA45_1C DEFAULT 
    LAYER Metal4 ;
        RECT -0.055000 -0.025000 0.055000 0.025000 ;
    LAYER Via4 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal5 ;
        RECT -0.025000 -0.055000 0.025000 0.055000 ;
END VIA45_1C

VIA VIA45_PG
    LAYER Metal4 ;
        RECT -0.200000 -0.050000 0.200000 0.050000 ;
    LAYER Via4 ;
        RECT -0.175000 -0.025000 -0.125000 0.025000 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
        RECT 0.125000 -0.025000 0.175000 0.025000 ;
    LAYER Metal5 ;
        RECT -0.200000 -0.050000 0.200000 0.050000 ;
END VIA45_PG

VIA VIA5_0_VH DEFAULT 
    LAYER Metal5 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
    LAYER Via5 ;
        RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal6 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
END VIA5_0_VH

VIA VIA56_PG
    LAYER Metal5 ;
        RECT -0.150000 -0.150000 0.150000 0.150000 ;
    LAYER Via5 ;
        RECT -0.150000 -0.150000 -0.100000 -0.100000 ;
        RECT -0.150000 0.100000 -0.100000 0.150000 ;
        RECT 0.100000 0.100000 0.150000 0.150000 ;
        RECT 0.100000 -0.150000 0.150000 -0.100000 ;
    LAYER Metal6 ;
        RECT -0.150000 -0.150000 0.150000 0.150000 ;
END VIA56_PG

VIA VIA6_0_HV DEFAULT 
    LAYER Metal6 ;
        RECT -0.065000 -0.035000 0.065000 0.035000 ;
    LAYER Via6 ;
        RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal7 ;
        RECT -0.035000 -0.065000 0.035000 0.065000 ;
END VIA6_0_HV

VIA VIA67_PG
    LAYER Metal6 ;
        RECT -0.170000 -0.170000 0.170000 0.170000 ;
    LAYER Via6 ;
        RECT -0.170000 -0.170000 -0.100000 -0.100000 ;
        RECT -0.170000 0.100000 -0.100000 0.170000 ;
        RECT 0.100000 0.100000 0.170000 0.170000 ;
        RECT 0.100000 -0.170000 0.170000 -0.100000 ;
    LAYER Metal7 ;
        RECT -0.170000 -0.170000 0.170000 0.170000 ;
END VIA67_PG

VIA VIA7_0_VH DEFAULT 
    LAYER Metal7 ;
        RECT -0.050000 -0.260000 0.050000 0.260000 ;
    LAYER Via7 ;
        RECT -0.050000 -0.050000 0.050000 0.050000 ;
    LAYER Metal8 ;
        RECT -0.260000 -0.050000 0.260000 0.050000 ;
END VIA7_0_VH

VIA VIA78_PG
    LAYER Metal7 ;
        RECT -0.170000 -0.170000 0.170000 0.170000 ;
    LAYER Via7 ;
        RECT -0.170000 -0.170000 -0.100000 -0.100000 ;
        RECT -0.170000 0.100000 -0.100000 0.170000 ;
        RECT 0.100000 0.100000 0.170000 0.170000 ;
        RECT 0.100000 -0.170000 0.170000 -0.100000 ;
    LAYER Metal8 ;
        RECT -0.170000 -0.170000 0.170000 0.170000 ;
END VIA78_PG

VIA VIA8_0_HV DEFAULT 
    LAYER Metal8 ;
        RECT -0.260000 -0.050000 0.260000 0.050000 ;
    LAYER Via8 ;
        RECT -0.050000 -0.050000 0.050000 0.050000 ;
    LAYER Metal9 ;
        RECT -0.050000 -0.260000 0.050000 0.260000 ;
END VIA8_0_HV

VIA VIA12_2C_W DEFAULT
    LAYER Metal1 ;
	RECT -0.150000 -0.055000 0.025000 0.055000 ;
    LAYER Via1 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
	RECT -0.150000 -0.025000 -0.100000 0.025000 ;
    LAYER Metal2 ;
	RECT -0.180000 -0.025000 0.055000 0.025000 ;
END VIA12_2C_W

VIA VIA12_2C_CH DEFAULT
    LAYER Metal1 ;
	RECT -0.087500 -0.055000 0.087500 0.055000 ;
    LAYER Via1 ;
	RECT 0.037500 -0.025000 0.087500 0.025000 ;
	RECT -0.087500 -0.025000 -0.037500 0.025000 ;
    LAYER Metal2 ;
	RECT -0.117500 -0.025000 0.117500 0.025000 ;
END VIA12_2C_CH

VIA VIA12_2C_E DEFAULT
    LAYER Metal1 ;
	RECT -0.025000 -0.055000 0.150000 0.055000 ;
    LAYER Via1 ;
	RECT 0.100000 -0.025000 0.150000 0.025000 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal2 ;
	RECT -0.055000 -0.025000 0.180000 0.025000 ;
END VIA12_2C_E

VIA VIA12_2C_S DEFAULT
    LAYER Metal1 ;
	RECT -0.025000 -0.180000 0.025000 0.055000 ;
    LAYER Via1 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
	RECT -0.025000 -0.150000 0.025000 -0.100000 ;
    LAYER Metal2 ;
	RECT -0.055000 -0.150000 0.055000 0.025000 ;
END VIA12_2C_S

VIA VIA12_2C_CV DEFAULT
    LAYER Metal1 ;
	RECT -0.025000 -0.117500 0.025000 0.117500 ;
    LAYER Via1 ;
	RECT -0.025000 0.037500 0.025000 0.087500 ;
	RECT -0.025000 -0.087500 0.025000 -0.037500 ;
    LAYER Metal2 ;
	RECT -0.055000 -0.087500 0.055000 0.087500 ;
END VIA12_2C_CV

VIA VIA12_2C_N DEFAULT
    LAYER Metal1 ;
	RECT -0.025000 -0.055000 0.025000 0.180000 ;
    LAYER Via1 ;
	RECT -0.025000 0.100000 0.025000 0.150000 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal2 ;
	RECT -0.055000 -0.025000 0.055000 0.150000 ;
END VIA12_2C_N

VIA VIA23_2C_W DEFAULT
    LAYER Metal2 ;
	RECT -0.180000 -0.025000 0.055000 0.025000 ;
    LAYER Via2 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
	RECT -0.150000 -0.025000 -0.100000 0.025000 ;
    LAYER Metal3 ;
	RECT -0.150000 -0.055000 0.025000 0.055000 ;
END VIA23_2C_W

VIA VIA23_2C_CH DEFAULT
    LAYER Metal2 ;
	RECT -0.117500 -0.025000 0.117500 0.025000 ;
    LAYER Via2 ;
	RECT 0.037500 -0.025000 0.087500 0.025000 ;
	RECT -0.087500 -0.025000 -0.037500 0.025000 ;
    LAYER Metal3 ;
	RECT -0.087500 -0.055000 0.087500 0.055000 ;
END VIA23_2C_CH

VIA VIA23_2C_E DEFAULT
    LAYER Metal2 ;
	RECT -0.055000 -0.025000 0.180000 0.025000 ;
    LAYER Via2 ;
	RECT 0.100000 -0.025000 0.150000 0.025000 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal3 ;
	RECT -0.025000 -0.055000 0.150000 0.055000 ;
END VIA23_2C_E

VIA VIA23_2C_S DEFAULT
    LAYER Metal2 ;
	RECT -0.055000 -0.150000 0.055000 0.025000 ;
    LAYER Via2 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
	RECT -0.025000 -0.150000 0.025000 -0.100000 ;
    LAYER Metal3 ;
	RECT -0.025000 -0.180000 0.025000 0.055000 ;
END VIA23_2C_S

VIA VIA23_2C_CV DEFAULT
    LAYER Metal2 ;
	RECT -0.055000 -0.087500 0.055000 0.087500 ;
    LAYER Via2 ;
	RECT -0.025000 0.037500 0.025000 0.087500 ;
	RECT -0.025000 -0.087500 0.025000 -0.037500 ;
    LAYER Metal3 ;
	RECT -0.025000 -0.117500 0.025000 0.117500 ;
END VIA23_2C_CV

VIA VIA23_2C_N DEFAULT
    LAYER Metal2 ;
	RECT -0.055000 -0.025000 0.055000 0.150000 ;
    LAYER Via2 ;
	RECT -0.025000 0.100000 0.025000 0.150000 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal3 ;
	RECT -0.025000 -0.055000 0.025000 0.180000 ;
END VIA23_2C_N

VIA VIA34_2C_W DEFAULT
    LAYER Metal3 ;
	RECT -0.150000 -0.055000 0.025000 0.055000 ;
    LAYER Via3 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
	RECT -0.150000 -0.025000 -0.100000 0.025000 ;
    LAYER Metal4 ;
	RECT -0.180000 -0.025000 0.055000 0.025000 ;
END VIA34_2C_W

VIA VIA34_2C_CH DEFAULT
    LAYER Metal3 ;
	RECT -0.087500 -0.055000 0.087500 0.055000 ;
    LAYER Via3 ;
	RECT 0.037500 -0.025000 0.087500 0.025000 ;
	RECT -0.087500 -0.025000 -0.037500 0.025000 ;
    LAYER Metal4 ;
	RECT -0.117500 -0.025000 0.117500 0.025000 ;
END VIA34_2C_CH

VIA VIA34_2C_E DEFAULT
    LAYER Metal3 ;
	RECT -0.025000 -0.055000 0.150000 0.055000 ;
    LAYER Via3 ;
	RECT 0.100000 -0.025000 0.150000 0.025000 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal4 ;
	RECT -0.055000 -0.025000 0.180000 0.025000 ;
END VIA34_2C_E

VIA VIA34_2C_S DEFAULT
    LAYER Metal3 ;
	RECT -0.025000 -0.180000 0.025000 0.055000 ;
    LAYER Via3 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
	RECT -0.025000 -0.150000 0.025000 -0.100000 ;
    LAYER Metal4 ;
	RECT -0.055000 -0.150000 0.055000 0.025000 ;
END VIA34_2C_S

VIA VIA34_2C_CV DEFAULT
    LAYER Metal3 ;
	RECT -0.025000 -0.117500 0.025000 0.117500 ;
    LAYER Via3 ;
	RECT -0.025000 0.037500 0.025000 0.087500 ;
	RECT -0.025000 -0.087500 0.025000 -0.037500 ;
    LAYER Metal4 ;
	RECT -0.055000 -0.087500 0.055000 0.087500 ;
END VIA34_2C_CV

VIA VIA34_2C_N DEFAULT
    LAYER Metal3 ;
	RECT -0.025000 -0.055000 0.025000 0.180000 ;
    LAYER Via3 ;
	RECT -0.025000 0.100000 0.025000 0.150000 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal4 ;
	RECT -0.055000 -0.025000 0.055000 0.150000 ;
END VIA34_2C_N

VIA VIA45_2C_W DEFAULT
    LAYER Metal4 ;
	RECT -0.180000 -0.025000 0.055000 0.025000 ;
    LAYER Via4 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
	RECT -0.150000 -0.025000 -0.100000 0.025000 ;
    LAYER Metal5 ;
	RECT -0.150000 -0.055000 0.025000 0.055000 ;
END VIA45_2C_W

VIA VIA45_2C_CH DEFAULT
    LAYER Metal4 ;
	RECT -0.117500 -0.025000 0.117500 0.025000 ;
    LAYER Via4 ;
	RECT 0.037500 -0.025000 0.087500 0.025000 ;
	RECT -0.087500 -0.025000 -0.037500 0.025000 ;
    LAYER Metal5 ;
	RECT -0.087500 -0.055000 0.087500 0.055000 ;
END VIA45_2C_CH

VIA VIA45_2C_E DEFAULT
    LAYER Metal4 ;
	RECT -0.055000 -0.025000 0.180000 0.025000 ;
    LAYER Via4 ;
	RECT 0.100000 -0.025000 0.150000 0.025000 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal5 ;
	RECT -0.025000 -0.055000 0.150000 0.055000 ;
END VIA45_2C_E

VIA VIA45_2C_S DEFAULT
    LAYER Metal4 ;
	RECT -0.055000 -0.150000 0.055000 0.025000 ;
    LAYER Via4 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
	RECT -0.025000 -0.150000 0.025000 -0.100000 ;
    LAYER Metal5 ;
	RECT -0.025000 -0.180000 0.025000 0.055000 ;
END VIA45_2C_S

VIA VIA45_2C_CV DEFAULT
    LAYER Metal4 ;
	RECT -0.055000 -0.087500 0.055000 0.087500 ;
    LAYER Via4 ;
	RECT -0.025000 0.037500 0.025000 0.087500 ;
	RECT -0.025000 -0.087500 0.025000 -0.037500 ;
    LAYER Metal5 ;
	RECT -0.025000 -0.117500 0.025000 0.117500 ;
END VIA45_2C_CV

VIA VIA45_2C_N DEFAULT
    LAYER Metal4 ;
	RECT -0.055000 -0.025000 0.055000 0.150000 ;
    LAYER Via4 ;
	RECT -0.025000 0.100000 0.025000 0.150000 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal5 ;
	RECT -0.025000 -0.055000 0.025000 0.180000 ;
END VIA45_2C_N

VIA VIA56_2C_W DEFAULT
    LAYER Metal5 ;
	RECT -0.150000 -0.055000 0.025000 0.055000 ;
    LAYER Via5 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
	RECT -0.150000 -0.025000 -0.100000 0.025000 ;
    LAYER Metal6 ;
	RECT -0.180000 -0.025000 0.055000 0.025000 ;
END VIA56_2C_W

VIA VIA56_2C_CH DEFAULT
    LAYER Metal5 ;
	RECT -0.087500 -0.055000 0.087500 0.055000 ;
    LAYER Via5 ;
	RECT 0.037500 -0.025000 0.087500 0.025000 ;
	RECT -0.087500 -0.025000 -0.037500 0.025000 ;
    LAYER Metal6 ;
	RECT -0.117500 -0.025000 0.117500 0.025000 ;
END VIA56_2C_CH

VIA VIA56_2C_E DEFAULT
    LAYER Metal5 ;
	RECT -0.025000 -0.055000 0.150000 0.055000 ;
    LAYER Via5 ;
	RECT 0.100000 -0.025000 0.150000 0.025000 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal6 ;
	RECT -0.055000 -0.025000 0.180000 0.025000 ;
END VIA56_2C_E

VIA VIA56_2C_S DEFAULT
    LAYER Metal5 ;
	RECT -0.025000 -0.180000 0.025000 0.055000 ;
    LAYER Via5 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
	RECT -0.025000 -0.150000 0.025000 -0.100000 ;
    LAYER Metal6 ;
	RECT -0.055000 -0.150000 0.055000 0.025000 ;
END VIA56_2C_S

VIA VIA56_2C_CV DEFAULT
    LAYER Metal5 ;
	RECT -0.025000 -0.117500 0.025000 0.117500 ;
    LAYER Via5 ;
	RECT -0.025000 0.037500 0.025000 0.087500 ;
	RECT -0.025000 -0.087500 0.025000 -0.037500 ;
    LAYER Metal6 ;
	RECT -0.055000 -0.087500 0.055000 0.087500 ;
END VIA56_2C_CV

VIA VIA56_2C_N DEFAULT
    LAYER Metal5 ;
	RECT -0.025000 -0.055000 0.025000 0.180000 ;
    LAYER Via5 ;
	RECT -0.025000 0.100000 0.025000 0.150000 ;
	RECT -0.025000 -0.025000 0.025000 0.025000 ;
    LAYER Metal6 ;
	RECT -0.055000 -0.025000 0.055000 0.150000 ;
END VIA56_2C_N

VIA VIA67_2C_W DEFAULT
    LAYER Metal6 ;
	RECT -0.235000 -0.035000 0.065000 0.035000 ;
    LAYER Via6 ;
	RECT -0.035000 -0.035000 0.035000 0.035000 ;
	RECT -0.205000 -0.035000 -0.135000 0.035000 ;
    LAYER Metal7 ;
	RECT -0.205000 -0.065000 0.035000 0.065000 ;
END VIA67_2C_W

VIA VIA67_2C_CH DEFAULT
    LAYER Metal6 ;
	RECT -0.150000 -0.035000 0.150000 0.035000 ;
    LAYER Via6 ;
	RECT 0.050000 -0.035000 0.120000 0.035000 ;
	RECT -0.120000 -0.035000 -0.050000 0.035000 ;
    LAYER Metal7 ;
	RECT -0.120000 -0.065000 0.120000 0.065000 ;
END VIA67_2C_CH

VIA VIA67_2C_E DEFAULT
    LAYER Metal6 ;
	RECT -0.065000 -0.035000 0.235000 0.035000 ;
    LAYER Via6 ;
	RECT 0.135000 -0.035000 0.205000 0.035000 ;
	RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal7 ;
	RECT -0.035000 -0.065000 0.205000 0.065000 ;
END VIA67_2C_E

VIA VIA67_2C_S DEFAULT
    LAYER Metal6 ;
	RECT -0.065000 -0.205000 0.065000 0.035000 ;
    LAYER Via6 ;
	RECT -0.035000 -0.035000 0.035000 0.035000 ;
	RECT -0.035000 -0.205000 0.035000 -0.135000 ;
    LAYER Metal7 ;
	RECT -0.035000 -0.235000 0.035000 0.065000 ;
END VIA67_2C_S

VIA VIA67_2C_CV DEFAULT
    LAYER Metal6 ;
	RECT -0.065000 -0.120000 0.065000 0.120000 ;
    LAYER Via6 ;
	RECT -0.035000 0.050000 0.035000 0.120000 ;
	RECT -0.035000 -0.120000 0.035000 -0.050000 ;
    LAYER Metal7 ;
	RECT -0.035000 -0.150000 0.035000 0.150000 ;
END VIA67_2C_CV

VIA VIA67_2C_N DEFAULT
    LAYER Metal6 ;
	RECT -0.065000 -0.035000 0.065000 0.205000 ;
    LAYER Via6 ;
	RECT -0.035000 0.135000 0.035000 0.205000 ;
	RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal7 ;
	RECT -0.035000 -0.065000 0.035000 0.235000 ;
END VIA67_2C_N

VIA VIA78_2C_W DEFAULT
    LAYER Metal7 ;
	RECT -0.205000 -0.065000 0.035000 0.065000 ;
    LAYER Via7 ;
	RECT -0.035000 -0.035000 0.035000 0.035000 ;
	RECT -0.205000 -0.035000 -0.135000 0.035000 ;
    LAYER Metal8 ;
	RECT -0.235000 -0.035000 0.065000 0.035000 ;
END VIA78_2C_W

VIA VIA78_2C_CH DEFAULT
    LAYER Metal7 ;
	RECT -0.120000 -0.065000 0.120000 0.065000 ;
    LAYER Via7 ;
	RECT 0.050000 -0.035000 0.120000 0.035000 ;
	RECT -0.120000 -0.035000 -0.050000 0.035000 ;
    LAYER Metal8 ;
	RECT -0.150000 -0.035000 0.150000 0.035000 ;
END VIA78_2C_CH

VIA VIA78_2C_E DEFAULT
    LAYER Metal7 ;
	RECT -0.035000 -0.065000 0.205000 0.065000 ;
    LAYER Via7 ;
	RECT 0.135000 -0.035000 0.205000 0.035000 ;
	RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal8 ;
	RECT -0.065000 -0.035000 0.235000 0.035000 ;
END VIA78_2C_E

VIA VIA78_2C_S DEFAULT
    LAYER Metal7 ;
	RECT -0.035000 -0.235000 0.035000 0.065000 ;
    LAYER Via7 ;
	RECT -0.035000 -0.035000 0.035000 0.035000 ;
	RECT -0.035000 -0.205000 0.035000 -0.135000 ;
    LAYER Metal8 ;
	RECT -0.065000 -0.205000 0.065000 0.035000 ;
END VIA78_2C_S

VIA VIA78_2C_CV DEFAULT
    LAYER Metal7 ;
	RECT -0.035000 -0.150000 0.035000 0.150000 ;
    LAYER Via7 ;
	RECT -0.035000 0.050000 0.035000 0.120000 ;
	RECT -0.035000 -0.120000 0.035000 -0.050000 ;
    LAYER Metal8 ;
	RECT -0.065000 -0.120000 0.065000 0.120000 ;
END VIA78_2C_CV

VIA VIA78_2C_N DEFAULT
    LAYER Metal7 ;
	RECT -0.035000 -0.065000 0.035000 0.235000 ;
    LAYER Via7 ;
	RECT -0.035000 0.135000 0.035000 0.205000 ;
	RECT -0.035000 -0.035000 0.035000 0.035000 ;
    LAYER Metal8 ;
	RECT -0.065000 -0.035000 0.065000 0.205000 ;
END VIA78_2C_N

VIARULE M4_M3 GENERATE DEFAULT
  LAYER Metal3 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER Via3 ;
    RECT -0.025 -0.025 0.025 0.025 ;
    SPACING 0.11 BY 0.11 ;
  LAYER Metal4 ;
    ENCLOSURE 0.005 0.03 ;
END M4_M3

VIARULE M5_M4 GENERATE DEFAULT
  LAYER Metal4 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER Via4 ;
    RECT -0.025 -0.025 0.025 0.025 ;
    SPACING 0.11 BY 0.11 ;
  LAYER Metal5 ;
    ENCLOSURE 0.005 0.03 ;
END M5_M4

VIARULE M6_M5 GENERATE DEFAULT
  LAYER Metal5 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER Via5 ;
    RECT -0.025 -0.025 0.025 0.025 ;
    SPACING 0.11 BY 0.11 ;
  LAYER Metal6 ;
    ENCLOSURE 0.005 0.03 ;
END M6_M5

VIARULE M7_M6 GENERATE DEFAULT
  LAYER Metal6 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER Via6 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.15 BY 0.15 ;
  LAYER Metal7 ;
    ENCLOSURE 0.005 0.03 ;
END M7_M6

VIARULE M8_M7 GENERATE DEFAULT
  LAYER Metal7 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER Via7 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.15 BY 0.15 ;
  LAYER Metal8 ;
    ENCLOSURE 0.005 0.03 ;
END M8_M7

SITE CoreSite
  CLASS CORE ;
  SIZE 0.1 BY 1.2 ;
END CoreSite

SITE pad
    SYMMETRY x y r90 ;
    CLASS pad ;
    SIZE 0.010 BY 23.5000 ;
END pad 

SITE corner
    SYMMETRY x y r90 ;
    CLASS pad ;
    SIZE 23.5000 BY 23.5000 ;
END corner


MACRO XNOR2X1
    CLASS CORE ;
    FOREIGN XNOR2X1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.400000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.440000 0.557000 0.542000 0.638000 ;
        RECT 0.440000 0.439000 0.501000 0.638000 ;
        RECT 0.162000 0.388000 0.223000 0.496000 ;
        RECT 0.407000 0.439000 0.501000 0.496000 ;
        RECT 0.162000 0.439000 0.232000 0.496000 ;
        RECT 0.162000 0.442000 0.501000 0.496000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.289000 0.555000 0.379000 0.636000 ;
        RECT 0.289000 0.555000 0.350000 0.761000 ;
        RECT 0.232000 0.706000 0.350000 0.761000 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.400000 1.280000 ;
        RECT 1.114000 1.078000 1.204000 1.280000 ;
        RECT 0.228000 1.078000 0.318000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.400000 0.080000 ;
        RECT 1.114000 -0.080000 1.204000 0.122000 ;
        RECT 0.235000 -0.080000 0.325000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.262000 0.707000 1.352000 0.788000 ;
        RECT 1.262000 0.279000 1.352000 0.360000 ;
        RECT 1.282000 0.573000 1.352000 0.788000 ;
        RECT 1.291000 0.279000 1.352000 0.788000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.040000 0.192000 0.138000 0.326000 ;
        RECT 0.040000 0.810000 0.138000 0.901000 ;
        RECT 0.973000 0.886000 1.063000 0.974000 ;
        RECT 1.140000 0.426000 1.229000 0.507000 ;
        RECT 0.927000 0.295000 1.035000 0.376000 ;
        RECT 0.774000 0.158000 0.864000 0.239000 ;
        RECT 0.477000 0.745000 0.664000 0.826000 ;
        RECT 0.477000 0.295000 0.567000 0.376000 ;
        RECT 1.140000 0.426000 1.201000 0.831000 ;
        RECT 0.974000 0.295000 1.035000 0.720000 ;
        RECT 0.725000 0.295000 0.786000 0.831000 ;
        RECT 0.603000 0.321000 0.664000 0.940000 ;
        RECT 0.455000 0.902000 0.516000 1.050000 ;
        RECT 0.386000 0.185000 0.447000 0.246000 ;
        RECT 0.077000 0.810000 0.138000 0.957000 ;
        RECT 0.040000 0.192000 0.101000 0.901000 ;
        RECT 0.912000 0.665000 1.035000 0.720000 ;
        RECT 0.725000 0.776000 1.201000 0.831000 ;
        RECT 0.477000 0.321000 0.664000 0.376000 ;
        RECT 0.455000 0.995000 0.719000 1.050000 ;
        RECT 0.077000 0.902000 0.516000 0.957000 ;
        RECT 0.603000 0.886000 1.063000 0.940000 ;
        RECT 0.386000 0.185000 0.864000 0.239000 ;
        RECT 0.040000 0.192000 0.447000 0.246000 ;
        RECT 0.077000 0.192000 0.101000 0.957000 ;
    END
END XNOR2X1

MACRO SDFFSHQX2
    CLASS CORE ;
    FOREIGN SDFFSHQX2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 4.900000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER Metal1 ;
        RECT 0.050000 0.906000 0.179000 1.008000 ;
        RECT 0.057000 0.906000 0.126000 1.027000 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.945000 0.435000 1.057000 0.557000 ;
        RECT 0.932000 0.439000 1.057000 0.494000 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 4.257000 0.679000 4.343000 0.761000 ;
        RECT 4.378000 0.281000 4.468000 0.362000 ;
        RECT 4.257000 0.679000 4.432000 0.760000 ;
        RECT 4.522000 0.307000 4.583000 0.733000 ;
        RECT 4.493000 0.307000 4.583000 0.367000 ;
        RECT 4.378000 0.307000 4.583000 0.362000 ;
        RECT 4.257000 0.679000 4.583000 0.733000 ;
        END
    END Q
    PIN SE
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.337000 0.485000 0.427000 0.565000 ;
        RECT 0.285000 0.485000 0.427000 0.552000 ;
        RECT 0.285000 0.444000 0.346000 0.552000 ;
        RECT 0.232000 0.439000 0.293000 0.499000 ;
        RECT 0.232000 0.444000 0.346000 0.499000 ;
        RECT 0.337000 0.444000 0.346000 0.565000 ;
        RECT 0.285000 0.439000 0.293000 0.552000 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.693000 0.548000 0.831000 0.657000 ;
        END
    END SI
    PIN SN
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 2.477000 0.870000 2.588000 0.973000 ;
        RECT 3.998000 0.518000 4.089000 0.599000 ;
        RECT 1.701000 0.581000 1.791000 0.662000 ;
        RECT 2.837000 0.870000 2.917000 0.973000 ;
        RECT 1.716000 0.573000 1.791000 0.662000 ;
        RECT 1.716000 0.573000 2.043000 0.639000 ;
        RECT 4.652000 0.502000 4.713000 0.894000 ;
        RECT 4.010000 0.518000 4.071000 0.894000 ;
        RECT 3.930000 0.839000 3.991000 1.025000 ;
        RECT 2.856000 0.870000 2.917000 1.025000 ;
        RECT 2.003000 0.585000 2.064000 1.039000 ;
        RECT 2.477000 0.870000 2.537000 1.039000 ;
        RECT 1.701000 0.581000 2.043000 0.639000 ;
        RECT 3.930000 0.839000 4.713000 0.894000 ;
        RECT 2.856000 0.970000 3.991000 1.025000 ;
        RECT 2.477000 0.870000 2.917000 0.925000 ;
        RECT 2.003000 0.985000 2.537000 1.039000 ;
        RECT 1.701000 0.585000 2.064000 0.639000 ;
        RECT 2.003000 0.573000 2.043000 1.039000 ;
        END
    END SN
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 1.727000 1.001000 1.942000 1.280000 ;
        RECT 0.000000 1.120000 4.900000 1.280000 ;
        RECT 4.459000 0.988000 4.549000 1.280000 ;
        RECT 4.061000 0.976000 4.151000 1.280000 ;
        RECT 2.665000 0.996000 2.755000 1.280000 ;
        RECT 0.805000 1.001000 0.895000 1.280000 ;
        RECT 0.199000 1.078000 0.289000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 4.900000 0.080000 ;
        RECT 0.742000 -0.080000 0.833000 0.122000 ;
        RECT 4.717000 -0.080000 4.807000 0.345000 ;
        RECT 3.740000 -0.080000 3.830000 0.122000 ;
        RECT 2.807000 -0.080000 2.897000 0.303000 ;
        RECT 1.635000 -0.080000 1.725000 0.214000 ;
        RECT 0.196000 -0.080000 0.286000 0.122000 ;
        RECT 2.439000 -0.080000 2.500000 0.311000 ;
        END
    END VSS
    OBS
        LAYER Metal1 ;
        RECT 3.374000 0.206000 3.477000 0.381000 ;
        RECT 3.183000 0.305000 3.273000 0.435000 ;
        RECT 2.001000 0.337000 2.091000 0.449000 ;
        RECT 3.731000 0.824000 3.821000 0.905000 ;
        RECT 3.712000 0.348000 3.802000 0.429000 ;
        RECT 3.655000 0.657000 3.745000 0.738000 ;
        RECT 3.633000 0.490000 3.723000 0.571000 ;
        RECT 2.992000 0.244000 3.082000 0.325000 ;
        RECT 2.866000 0.733000 2.956000 0.814000 ;
        RECT 2.616000 0.265000 2.706000 0.346000 ;
        RECT 2.475000 0.733000 2.565000 0.814000 ;
        RECT 2.160000 0.848000 2.250000 0.929000 ;
        RECT 1.937000 0.171000 2.027000 0.252000 ;
        RECT 1.808000 0.779000 1.898000 0.860000 ;
        RECT 1.522000 0.517000 1.612000 0.598000 ;
        RECT 1.399000 0.930000 1.489000 1.011000 ;
        RECT 1.157000 0.442000 1.248000 0.523000 ;
        RECT 0.408000 0.343000 0.593000 0.424000 ;
        RECT 0.382000 0.150000 0.472000 0.231000 ;
        RECT 0.048000 0.746000 0.138000 0.827000 ;
        RECT 0.048000 0.323000 0.138000 0.404000 ;
        RECT 2.305000 0.835000 2.414000 0.915000 ;
        RECT 3.633000 0.490000 3.788000 0.561000 ;
        RECT 3.731000 0.824000 3.869000 0.892000 ;
        RECT 0.038000 0.746000 0.138000 0.814000 ;
        RECT 2.160000 0.848000 2.414000 0.915000 ;
        RECT 0.526000 0.315000 0.593000 0.424000 ;
        RECT 4.152000 0.206000 4.213000 0.554000 ;
        RECT 3.808000 0.506000 3.869000 0.892000 ;
        RECT 3.727000 0.348000 3.788000 0.561000 ;
        RECT 3.416000 0.206000 3.477000 0.915000 ;
        RECT 3.374000 0.189000 3.435000 0.381000 ;
        RECT 3.226000 0.380000 3.287000 0.801000 ;
        RECT 3.021000 0.189000 3.082000 0.325000 ;
        RECT 2.645000 0.265000 2.706000 0.435000 ;
        RECT 2.353000 0.417000 2.414000 0.915000 ;
        RECT 2.254000 0.336000 2.315000 0.471000 ;
        RECT 2.227000 0.161000 2.288000 0.390000 ;
        RECT 2.225000 0.533000 2.286000 0.685000 ;
        RECT 2.129000 0.446000 2.190000 0.588000 ;
        RECT 2.030000 0.337000 2.091000 0.501000 ;
        RECT 1.844000 0.198000 1.905000 0.338000 ;
        RECT 1.537000 0.394000 1.598000 0.846000 ;
        RECT 1.323000 0.283000 1.384000 0.850000 ;
        RECT 1.201000 0.732000 1.262000 0.998000 ;
        RECT 1.172000 0.442000 1.233000 0.787000 ;
        RECT 1.112000 0.156000 1.173000 0.261000 ;
        RECT 1.079000 0.856000 1.140000 0.979000 ;
        RECT 0.668000 0.856000 0.729000 1.023000 ;
        RECT 0.534000 0.732000 0.595000 0.913000 ;
        RECT 0.532000 0.315000 0.593000 0.677000 ;
        RECT 0.412000 0.623000 0.473000 0.779000 ;
        RECT 0.411000 0.150000 0.472000 0.261000 ;
        RECT 0.289000 0.773000 0.350000 0.913000 ;
        RECT 0.038000 0.349000 0.099000 0.814000 ;
        RECT 4.152000 0.499000 4.429000 0.554000 ;
        RECT 3.727000 0.506000 3.869000 0.561000 ;
        RECT 3.633000 0.670000 3.745000 0.725000 ;
        RECT 3.633000 0.506000 3.802000 0.561000 ;
        RECT 3.477000 0.670000 3.655000 0.725000 ;
        RECT 3.477000 0.206000 4.213000 0.261000 ;
        RECT 3.416000 0.670000 3.633000 0.725000 ;
        RECT 3.374000 0.206000 3.869000 0.261000 ;
        RECT 3.021000 0.189000 3.435000 0.244000 ;
        RECT 2.645000 0.380000 3.287000 0.435000 ;
        RECT 2.475000 0.746000 3.354000 0.801000 ;
        RECT 2.353000 0.489000 3.162000 0.544000 ;
        RECT 2.129000 0.533000 2.286000 0.588000 ;
        RECT 2.030000 0.446000 2.190000 0.501000 ;
        RECT 1.537000 0.394000 2.091000 0.449000 ;
        RECT 1.323000 0.283000 1.905000 0.338000 ;
        RECT 1.201000 0.943000 1.489000 0.998000 ;
        RECT 1.112000 0.156000 1.209000 0.211000 ;
        RECT 0.668000 0.856000 1.140000 0.911000 ;
        RECT 0.534000 0.732000 1.262000 0.787000 ;
        RECT 0.526000 0.315000 0.920000 0.370000 ;
        RECT 0.443000 0.968000 0.729000 1.023000 ;
        RECT 0.411000 0.206000 1.173000 0.261000 ;
        RECT 0.289000 0.858000 0.595000 0.913000 ;
        RECT 0.038000 0.349000 0.138000 0.404000 ;
        RECT 3.057000 0.861000 3.477000 0.915000 ;
        RECT 2.254000 0.417000 2.414000 0.471000 ;
        RECT 2.227000 0.336000 2.315000 0.390000 ;
        RECT 2.117000 0.161000 2.288000 0.215000 ;
        RECT 1.844000 0.198000 2.027000 0.252000 ;
        RECT 1.537000 0.792000 1.898000 0.846000 ;
        RECT 1.267000 0.323000 1.384000 0.377000 ;
        RECT 0.412000 0.623000 0.593000 0.677000 ;
        RECT 0.048000 0.773000 0.350000 0.827000 ;
        RECT 0.048000 0.323000 0.099000 0.827000 ;
        RECT 3.226000 0.305000 3.273000 0.801000 ;
        RECT 2.254000 0.161000 2.288000 0.471000 ;
        RECT 1.201000 0.442000 1.233000 0.998000 ;
        RECT 3.416000 0.189000 3.435000 0.915000 ;
        RECT 3.808000 0.506000 3.821000 0.905000 ;
    END
END SDFFSHQX2

MACRO SDFFSHQX1
    CLASS CORE ;
    FOREIGN SDFFSHQX1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 4.200000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER Metal1 ;
        RECT 0.208000 0.439000 0.273000 0.565000 ;
        RECT 0.208000 0.439000 0.269000 0.567000 ;
        RECT 0.160000 0.511000 0.221000 0.598000 ;
        RECT 0.160000 0.511000 0.269000 0.567000 ;
        RECT 0.208000 0.439000 0.293000 0.494000 ;
        RECT 0.160000 0.511000 0.273000 0.565000 ;
        RECT 0.208000 0.439000 0.221000 0.598000 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.031000 0.421000 1.172000 0.536000 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 4.028000 0.204000 4.143000 0.290000 ;
        RECT 4.062000 0.627000 4.143000 0.715000 ;
        RECT 4.062000 0.204000 4.143000 0.307000 ;
        RECT 3.745000 0.738000 3.835000 0.819000 ;
        RECT 4.082000 0.204000 4.143000 0.715000 ;
        RECT 3.774000 0.661000 3.835000 0.819000 ;
        RECT 3.774000 0.661000 4.143000 0.715000 ;
        END
    END Q
    PIN SE
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.374000 0.539000 0.496000 0.669000 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.737000 0.344000 0.818000 0.439000 ;
        RECT 0.720000 0.593000 0.810000 0.674000 ;
        RECT 0.703000 0.331000 0.793000 0.412000 ;
        RECT 0.720000 0.593000 0.818000 0.661000 ;
        RECT 0.703000 0.344000 0.818000 0.412000 ;
        RECT 0.757000 0.344000 0.818000 0.661000 ;
        RECT 0.737000 0.331000 0.793000 0.439000 ;
        RECT 0.757000 0.344000 0.810000 0.674000 ;
        RECT 0.757000 0.331000 0.793000 0.674000 ;
        END
    END SI
    PIN SN
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.804000 0.608000 2.043000 0.701000 ;
        RECT 3.607000 0.502000 3.698000 0.583000 ;
        RECT 1.804000 0.633000 2.136000 0.701000 ;
        RECT 3.732000 0.439000 3.793000 0.500000 ;
        RECT 3.637000 0.445000 3.698000 0.583000 ;
        RECT 3.517000 0.529000 3.578000 0.994000 ;
        RECT 2.075000 0.633000 2.136000 0.994000 ;
        RECT 1.982000 0.573000 2.043000 0.701000 ;
        RECT 3.637000 0.445000 3.793000 0.500000 ;
        RECT 2.075000 0.939000 3.578000 0.994000 ;
        RECT 3.517000 0.529000 3.698000 0.583000 ;
        END
    END SN
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 1.763000 1.001000 2.013000 1.280000 ;
        RECT 0.000000 1.120000 4.200000 1.280000 ;
        RECT 2.369000 1.078000 2.466000 1.280000 ;
        RECT 3.936000 0.805000 4.026000 1.280000 ;
        RECT 3.590000 1.078000 3.680000 1.280000 ;
        RECT 3.218000 1.078000 3.308000 1.280000 ;
        RECT 0.202000 1.078000 0.292000 1.280000 ;
        RECT 0.925000 1.002000 0.986000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 4.200000 0.080000 ;
        RECT 3.663000 -0.080000 3.753000 0.122000 ;
        RECT 3.222000 -0.080000 3.312000 0.122000 ;
        RECT 1.681000 -0.080000 1.771000 0.186000 ;
        RECT 0.745000 -0.080000 0.835000 0.122000 ;
        RECT 0.196000 -0.080000 0.286000 0.206000 ;
        RECT 2.459000 -0.080000 2.520000 0.290000 ;
        END
    END VSS
    OBS
        LAYER Metal1 ;
        RECT 2.040000 0.318000 2.141000 0.475000 ;
        RECT 3.903000 0.502000 3.993000 0.583000 ;
        RECT 3.387000 0.165000 3.481000 0.246000 ;
        RECT 3.077000 0.629000 3.167000 0.710000 ;
        RECT 2.636000 0.257000 2.726000 0.338000 ;
        RECT 2.233000 0.295000 2.323000 0.376000 ;
        RECT 2.197000 0.790000 2.287000 0.871000 ;
        RECT 2.158000 0.150000 2.248000 0.231000 ;
        RECT 1.953000 0.171000 2.043000 0.252000 ;
        RECT 1.845000 0.795000 1.936000 0.876000 ;
        RECT 1.579000 0.426000 1.743000 0.507000 ;
        RECT 1.409000 0.700000 1.499000 0.781000 ;
        RECT 1.335000 0.862000 1.425000 0.943000 ;
        RECT 1.319000 0.190000 1.409000 0.271000 ;
        RECT 1.250000 0.438000 1.340000 0.519000 ;
        RECT 1.123000 0.825000 1.213000 0.906000 ;
        RECT 1.106000 0.257000 1.196000 0.338000 ;
        RECT 0.445000 0.346000 0.536000 0.427000 ;
        RECT 0.048000 0.743000 0.138000 0.824000 ;
        RECT 0.037000 0.331000 0.138000 0.412000 ;
        RECT 1.106000 0.206000 1.183000 0.338000 ;
        RECT 0.460000 0.346000 0.536000 0.444000 ;
        RECT 2.390000 0.804000 2.483000 0.874000 ;
        RECT 2.158000 0.163000 2.294000 0.231000 ;
        RECT 2.197000 0.804000 2.483000 0.871000 ;
        RECT 1.319000 0.204000 1.493000 0.271000 ;
        RECT 0.037000 0.743000 0.138000 0.807000 ;
        RECT 2.935000 0.192000 2.998000 0.290000 ;
        RECT 1.430000 0.204000 1.493000 0.325000 ;
        RECT 3.903000 0.306000 3.964000 0.583000 ;
        RECT 3.451000 0.192000 3.512000 0.361000 ;
        RECT 3.393000 0.629000 3.454000 0.750000 ;
        RECT 3.328000 0.314000 3.389000 0.683000 ;
        RECT 3.126000 0.192000 3.187000 0.539000 ;
        RECT 2.911000 0.485000 2.972000 0.760000 ;
        RECT 2.787000 0.345000 2.848000 0.582000 ;
        RECT 2.683000 0.527000 2.744000 0.614000 ;
        RECT 2.636000 0.257000 2.697000 0.437000 ;
        RECT 2.557000 0.382000 2.618000 0.760000 ;
        RECT 2.422000 0.380000 2.483000 0.874000 ;
        RECT 2.335000 0.321000 2.396000 0.435000 ;
        RECT 2.233000 0.163000 2.294000 0.376000 ;
        RECT 2.213000 0.431000 2.274000 0.615000 ;
        RECT 2.080000 0.318000 2.141000 0.486000 ;
        RECT 1.865000 0.198000 1.926000 0.325000 ;
        RECT 1.682000 0.420000 1.743000 0.850000 ;
        RECT 1.560000 0.563000 1.621000 0.917000 ;
        RECT 1.430000 0.204000 1.491000 0.618000 ;
        RECT 1.265000 0.438000 1.326000 0.755000 ;
        RECT 0.917000 0.601000 0.978000 0.787000 ;
        RECT 0.802000 0.851000 0.863000 1.025000 ;
        RECT 0.679000 0.732000 0.740000 0.915000 ;
        RECT 0.557000 0.389000 0.618000 0.789000 ;
        RECT 0.396000 0.152000 0.457000 0.261000 ;
        RECT 0.077000 0.743000 0.138000 0.915000 ;
        RECT 0.037000 0.331000 0.098000 0.807000 ;
        RECT 3.451000 0.306000 3.964000 0.361000 ;
        RECT 2.800000 0.705000 2.972000 0.760000 ;
        RECT 2.787000 0.345000 3.060000 0.400000 ;
        RECT 2.683000 0.527000 2.848000 0.582000 ;
        RECT 2.557000 0.705000 2.677000 0.760000 ;
        RECT 2.557000 0.382000 2.697000 0.437000 ;
        RECT 2.390000 0.819000 3.051000 0.874000 ;
        RECT 2.335000 0.380000 2.483000 0.435000 ;
        RECT 2.233000 0.321000 2.396000 0.376000 ;
        RECT 2.080000 0.431000 2.274000 0.486000 ;
        RECT 1.682000 0.795000 1.936000 0.850000 ;
        RECT 1.682000 0.420000 2.141000 0.475000 ;
        RECT 1.430000 0.563000 1.621000 0.618000 ;
        RECT 1.430000 0.270000 1.926000 0.325000 ;
        RECT 1.335000 0.862000 1.621000 0.917000 ;
        RECT 1.265000 0.700000 1.499000 0.755000 ;
        RECT 0.917000 0.601000 1.326000 0.656000 ;
        RECT 0.802000 0.851000 1.213000 0.906000 ;
        RECT 0.679000 0.732000 0.978000 0.787000 ;
        RECT 0.460000 0.389000 0.618000 0.444000 ;
        RECT 0.438000 0.970000 0.863000 1.025000 ;
        RECT 0.396000 0.206000 1.183000 0.261000 ;
        RECT 3.077000 0.629000 3.454000 0.683000 ;
        RECT 2.935000 0.192000 3.512000 0.246000 ;
        RECT 2.911000 0.485000 3.187000 0.539000 ;
        RECT 2.828000 0.236000 2.998000 0.290000 ;
        RECT 2.213000 0.561000 2.360000 0.615000 ;
        RECT 1.865000 0.198000 2.043000 0.252000 ;
        RECT 0.404000 0.735000 0.618000 0.789000 ;
        RECT 0.077000 0.861000 0.740000 0.915000 ;
        RECT 2.197000 0.819000 3.051000 0.871000 ;
        RECT 0.048000 0.331000 0.098000 0.824000 ;
        RECT 3.451000 0.165000 3.481000 0.361000 ;
        RECT 0.077000 0.331000 0.098000 0.915000 ;
        RECT 2.233000 0.150000 2.248000 0.376000 ;
    END
END SDFFSHQX1

MACRO SDFFRHQX4
    CLASS CORE ;
    FOREIGN SDFFRHQX4 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 6.400000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER Metal1 ;
        RECT 0.165000 0.476000 0.290000 0.627000 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.044000 0.706000 1.206000 0.792000 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 6.091000 0.349000 6.190000 0.767000 ;
        RECT 6.244000 0.707000 6.333000 0.931000 ;
        RECT 5.918000 0.179000 6.007000 0.404000 ;
        RECT 5.573000 0.707000 5.662000 0.931000 ;
        RECT 5.540000 0.179000 5.629000 0.402000 ;
        RECT 6.244000 0.706000 6.319000 0.931000 ;
        RECT 5.555000 0.179000 5.629000 0.404000 ;
        RECT 6.091000 0.706000 6.319000 0.767000 ;
        RECT 6.091000 0.707000 6.333000 0.767000 ;
        RECT 5.573000 0.712000 6.333000 0.767000 ;
        RECT 5.555000 0.349000 6.190000 0.404000 ;
        RECT 5.540000 0.349000 6.190000 0.402000 ;
        END
    END Q
    PIN RN
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 4.529000 0.437000 4.787000 0.500000 ;
        RECT 4.527000 0.437000 4.787000 0.492000 ;
        END
    END RN
    PIN SE
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.921000 0.562000 0.981000 0.627000 ;
        RECT 0.769000 0.454000 0.829000 0.617000 ;
        RECT 0.769000 0.562000 1.090000 0.617000 ;
        RECT 0.689000 0.454000 0.829000 0.508000 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.729000 0.671000 0.828000 0.806000 ;
        END
    END SI
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 6.400000 1.280000 ;
        RECT 1.783000 1.078000 1.873000 1.280000 ;
        RECT 5.909000 0.910000 5.998000 1.280000 ;
        RECT 4.792000 1.078000 4.881000 1.280000 ;
        RECT 4.361000 0.989000 4.450000 1.280000 ;
        RECT 3.052000 1.078000 3.141000 1.280000 ;
        RECT 2.279000 1.078000 2.368000 1.280000 ;
        RECT 0.257000 1.078000 0.346000 1.280000 ;
        RECT 5.252000 0.742000 5.312000 1.280000 ;
        RECT 2.681000 0.982000 2.741000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 6.400000 0.080000 ;
        RECT 6.106000 -0.080000 6.196000 0.235000 ;
        RECT 1.804000 -0.080000 1.894000 0.216000 ;
        RECT 5.729000 -0.080000 5.818000 0.235000 ;
        RECT 4.834000 -0.080000 4.923000 0.122000 ;
        RECT 4.446000 -0.080000 4.535000 0.268000 ;
        RECT 2.994000 -0.080000 3.083000 0.299000 ;
        RECT 2.617000 -0.080000 2.706000 0.340000 ;
        RECT 0.962000 -0.080000 1.051000 0.122000 ;
        RECT 0.248000 -0.080000 0.337000 0.122000 ;
        RECT 5.316000 -0.080000 5.377000 0.360000 ;
        RECT 2.207000 -0.080000 2.267000 0.366000 ;
        RECT 2.192000 0.315000 2.281000 0.366000 ;
        END
    END VSS
    OBS
        LAYER Metal1 ;
        RECT 3.469000 0.285000 3.613000 0.458000 ;
        RECT 2.053000 0.699000 2.443000 0.792000 ;
        RECT 1.900000 0.480000 1.993000 0.615000 ;
        RECT 0.043000 0.729000 0.136000 0.952000 ;
        RECT 0.043000 0.167000 0.136000 0.360000 ;
        RECT 3.712000 0.161000 3.801000 0.329000 ;
        RECT 5.196000 0.506000 5.314000 0.594000 ;
        RECT 2.018000 0.294000 2.116000 0.381000 ;
        RECT 1.001000 0.344000 1.090000 0.431000 ;
        RECT 1.512000 0.480000 1.616000 0.563000 ;
        RECT 4.635000 0.236000 4.724000 0.317000 ;
        RECT 4.083000 0.262000 4.179000 0.343000 ;
        RECT 2.806000 0.270000 2.895000 0.351000 ;
        RECT 2.650000 0.655000 2.739000 0.736000 ;
        RECT 1.924000 0.698000 2.116000 0.779000 ;
        RECT 1.726000 0.612000 1.815000 0.693000 ;
        RECT 1.549000 0.650000 1.638000 0.731000 ;
        RECT 1.498000 0.214000 1.587000 0.295000 ;
        RECT 0.455000 0.476000 0.544000 0.557000 ;
        RECT 0.605000 0.208000 0.695000 0.287000 ;
        RECT 4.010000 0.627000 4.143000 0.704000 ;
        RECT 4.649000 0.192000 4.724000 0.317000 ;
        RECT 3.474000 0.692000 3.549000 0.792000 ;
        RECT 1.309000 0.208000 1.401000 0.275000 ;
        RECT 2.053000 0.698000 2.116000 0.792000 ;
        RECT 4.231000 0.862000 4.292000 1.039000 ;
        RECT 3.488000 0.285000 3.549000 0.792000 ;
        RECT 3.353000 0.815000 3.414000 0.915000 ;
        RECT 3.336000 0.421000 3.397000 0.580000 ;
        RECT 3.201000 0.954000 3.262000 1.039000 ;
        RECT 3.197000 0.285000 3.258000 0.425000 ;
        RECT 2.834000 0.270000 2.895000 0.425000 ;
        RECT 2.247000 0.919000 2.308000 0.994000 ;
        RECT 1.563000 0.650000 1.624000 0.994000 ;
        RECT 1.424000 0.508000 1.485000 0.818000 ;
        RECT 1.386000 0.350000 1.447000 0.437000 ;
        RECT 0.043000 0.167000 0.104000 0.952000 ;
        RECT 5.196000 0.192000 5.256000 0.594000 ;
        RECT 5.132000 0.539000 5.192000 0.994000 ;
        RECT 5.075000 0.301000 5.135000 0.423000 ;
        RECT 5.011000 0.524000 5.071000 0.885000 ;
        RECT 4.884000 0.368000 4.944000 0.775000 ;
        RECT 4.647000 0.751000 4.707000 0.885000 ;
        RECT 4.513000 0.862000 4.573000 0.994000 ;
        RECT 4.407000 0.524000 4.467000 0.665000 ;
        RECT 4.285000 0.649000 4.345000 0.806000 ;
        RECT 4.111000 0.762000 4.171000 0.915000 ;
        RECT 4.083000 0.161000 4.143000 0.704000 ;
        RECT 3.863000 0.285000 3.923000 0.458000 ;
        RECT 3.626000 0.600000 3.686000 0.682000 ;
        RECT 3.057000 0.660000 3.117000 0.746000 ;
        RECT 2.922000 0.525000 2.982000 0.870000 ;
        RECT 2.802000 0.808000 2.862000 1.008000 ;
        RECT 2.664000 0.423000 2.724000 0.736000 ;
        RECT 2.542000 0.919000 2.602000 1.005000 ;
        RECT 2.504000 0.546000 2.564000 0.863000 ;
        RECT 2.456000 0.300000 2.516000 0.477000 ;
        RECT 2.427000 0.161000 2.487000 0.381000 ;
        RECT 2.056000 0.294000 2.116000 0.792000 ;
        RECT 1.755000 0.612000 1.815000 0.752000 ;
        RECT 1.512000 0.214000 1.572000 0.563000 ;
        RECT 1.266000 0.382000 1.326000 0.932000 ;
        RECT 0.607000 0.775000 0.667000 0.932000 ;
        RECT 0.485000 0.885000 0.545000 1.042000 ;
        RECT 0.469000 0.256000 0.529000 0.720000 ;
        RECT 1.266000 0.874000 1.624000 0.932000 ;
        RECT 5.196000 0.506000 5.902000 0.561000 ;
        RECT 5.132000 0.539000 5.314000 0.594000 ;
        RECT 4.884000 0.368000 5.135000 0.423000 ;
        RECT 4.647000 0.830000 5.071000 0.885000 ;
        RECT 4.513000 0.939000 5.192000 0.994000 ;
        RECT 4.285000 0.751000 4.707000 0.806000 ;
        RECT 4.252000 0.524000 4.467000 0.579000 ;
        RECT 4.231000 0.862000 4.573000 0.917000 ;
        RECT 4.010000 0.649000 4.345000 0.704000 ;
        RECT 3.626000 0.627000 4.143000 0.682000 ;
        RECT 3.474000 0.737000 3.900000 0.792000 ;
        RECT 2.922000 0.815000 3.414000 0.870000 ;
        RECT 2.834000 0.370000 3.258000 0.425000 ;
        RECT 2.664000 0.525000 3.397000 0.580000 ;
        RECT 2.504000 0.808000 2.862000 0.863000 ;
        RECT 2.247000 0.919000 2.602000 0.974000 ;
        RECT 2.177000 0.546000 2.564000 0.601000 ;
        RECT 1.563000 0.939000 2.308000 0.994000 ;
        RECT 1.512000 0.480000 1.993000 0.535000 ;
        RECT 1.424000 0.508000 1.616000 0.563000 ;
        RECT 1.266000 0.382000 1.447000 0.437000 ;
        RECT 0.607000 0.877000 1.624000 0.932000 ;
        RECT 0.605000 0.208000 1.401000 0.263000 ;
        RECT 0.485000 0.987000 1.300000 1.042000 ;
        RECT 0.469000 0.344000 1.090000 0.399000 ;
        RECT 0.440000 0.665000 0.529000 0.720000 ;
        RECT 0.422000 0.256000 0.529000 0.311000 ;
        RECT 0.043000 0.775000 0.667000 0.830000 ;
        RECT 4.649000 0.192000 5.256000 0.246000 ;
        RECT 4.407000 0.611000 4.944000 0.665000 ;
        RECT 3.863000 0.285000 3.990000 0.339000 ;
        RECT 3.469000 0.404000 3.923000 0.458000 ;
        RECT 3.353000 0.861000 4.171000 0.915000 ;
        RECT 3.324000 0.161000 4.143000 0.215000 ;
        RECT 3.201000 0.985000 4.292000 1.039000 ;
        RECT 3.197000 0.285000 3.613000 0.339000 ;
        RECT 3.057000 0.692000 3.549000 0.746000 ;
        RECT 2.802000 0.954000 3.262000 1.008000 ;
        RECT 2.456000 0.423000 2.724000 0.477000 ;
        RECT 2.331000 0.161000 2.487000 0.215000 ;
        RECT 1.755000 0.698000 2.116000 0.752000 ;
        RECT 0.451000 0.885000 0.545000 0.939000 ;
        RECT 2.456000 0.161000 2.487000 0.477000 ;
    END
END SDFFRHQX4

MACRO SDFFRHQX1
    CLASS CORE ;
    FOREIGN SDFFRHQX1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 4.400000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER Metal1 ;
        RECT 0.168000 0.517000 0.295000 0.627000 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.035000 0.417000 1.195000 0.502000 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 4.248000 0.829000 4.355000 0.973000 ;
        RECT 4.248000 0.829000 4.339000 1.021000 ;
        RECT 3.965000 0.174000 4.056000 0.255000 ;
        RECT 4.281000 0.706000 4.355000 0.973000 ;
        RECT 4.295000 0.296000 4.356000 0.761000 ;
        RECT 3.995000 0.174000 4.056000 0.351000 ;
        RECT 4.295000 0.296000 4.355000 0.973000 ;
        RECT 4.281000 0.706000 4.339000 1.021000 ;
        RECT 4.281000 0.706000 4.356000 0.761000 ;
        RECT 3.995000 0.296000 4.356000 0.351000 ;
        RECT 4.295000 0.296000 4.339000 1.021000 ;
        END
    END Q
    PIN RN
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 3.800000 0.693000 4.011000 0.776000 ;
        END
    END RN
    PIN SE
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.380000 0.348000 0.492000 0.543000 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.787000 0.488000 0.877000 0.569000 ;
        RECT 0.801000 0.488000 0.877000 0.627000 ;
        RECT 0.801000 0.567000 0.999000 0.627000 ;
        END
    END SI
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 4.400000 1.280000 ;
        RECT 3.284000 1.078000 3.395000 1.280000 ;
        RECT 2.517000 1.078000 2.628000 1.280000 ;
        RECT 3.907000 0.857000 3.997000 1.280000 ;
        RECT 1.691000 0.963000 1.781000 1.280000 ;
        RECT 0.843000 1.001000 0.933000 1.280000 ;
        RECT 0.155000 0.932000 0.245000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 3.601000 -0.080000 3.852000 0.122000 ;
        RECT 0.000000 -0.080000 4.400000 0.080000 ;
        RECT 4.157000 -0.080000 4.248000 0.211000 ;
        RECT 2.425000 -0.080000 2.516000 0.254000 ;
        RECT 1.685000 -0.080000 1.776000 0.327000 ;
        RECT 0.197000 -0.080000 0.288000 0.122000 ;
        RECT 3.207000 -0.080000 3.297000 0.122000 ;
        RECT 0.747000 -0.080000 0.837000 0.122000 ;
        END
    END VSS
    OBS
        LAYER Metal1 ;
        RECT 3.527000 0.526000 3.679000 0.638000 ;
        RECT 2.596000 0.548000 2.720000 0.644000 ;
        RECT 3.269000 0.614000 3.360000 0.833000 ;
        RECT 0.384000 0.152000 0.475000 0.261000 ;
        RECT 1.109000 0.206000 1.200000 0.293000 ;
        RECT 0.821000 0.317000 0.911000 0.402000 ;
        RECT 4.093000 0.407000 4.184000 0.488000 ;
        RECT 3.713000 0.952000 3.804000 1.033000 ;
        RECT 3.601000 0.327000 3.692000 0.408000 ;
        RECT 3.388000 0.336000 3.479000 0.417000 ;
        RECT 3.211000 0.614000 3.360000 0.695000 ;
        RECT 2.927000 0.382000 3.017000 0.463000 ;
        RECT 2.925000 0.802000 3.016000 0.883000 ;
        RECT 2.843000 0.223000 2.933000 0.304000 ;
        RECT 2.733000 0.802000 2.843000 0.883000 ;
        RECT 2.629000 0.240000 2.720000 0.321000 ;
        RECT 2.381000 0.798000 2.472000 0.879000 ;
        RECT 2.287000 0.364000 2.384000 0.445000 ;
        RECT 2.123000 0.614000 2.213000 0.695000 ;
        RECT 1.880000 0.795000 1.987000 0.876000 ;
        RECT 1.859000 0.398000 1.949000 0.479000 ;
        RECT 1.581000 0.483000 1.672000 0.564000 ;
        RECT 1.459000 0.890000 1.549000 0.971000 ;
        RECT 1.323000 0.223000 1.413000 0.304000 ;
        RECT 0.821000 0.317000 0.912000 0.398000 ;
        RECT 0.600000 0.595000 0.691000 0.676000 ;
        RECT 0.557000 0.348000 0.649000 0.429000 ;
        RECT 0.533000 0.938000 0.624000 1.019000 ;
        RECT 0.400000 0.667000 0.491000 0.748000 ;
        RECT 0.044000 0.688000 0.139000 0.769000 ;
        RECT 0.044000 0.317000 0.139000 0.398000 ;
        RECT 0.572000 0.348000 0.649000 0.663000 ;
        RECT 2.857000 0.206000 2.933000 0.304000 ;
        RECT 3.497000 0.952000 3.804000 1.020000 ;
        RECT 2.904000 0.395000 3.017000 0.463000 ;
        RECT 2.123000 0.627000 2.247000 0.695000 ;
        RECT 1.859000 0.411000 1.987000 0.479000 ;
        RECT 0.572000 0.595000 0.691000 0.663000 ;
        RECT 3.295000 0.206000 3.393000 0.273000 ;
        RECT 3.497000 0.573000 3.679000 0.638000 ;
        RECT 3.617000 0.327000 3.679000 0.638000 ;
        RECT 3.497000 0.573000 3.559000 1.020000 ;
        RECT 2.781000 0.380000 2.843000 0.883000 ;
        RECT 2.473000 0.501000 2.535000 0.694000 ;
        RECT 2.185000 0.627000 2.247000 0.994000 ;
        RECT 1.925000 0.411000 1.987000 0.876000 ;
        RECT 1.257000 0.436000 1.319000 0.945000 ;
        RECT 0.429000 0.608000 0.491000 0.748000 ;
        RECT 0.077000 0.688000 0.139000 0.860000 ;
        RECT 3.779000 0.206000 3.840000 0.462000 ;
        RECT 3.299000 0.362000 3.360000 0.833000 ;
        RECT 3.080000 0.206000 3.141000 0.857000 ;
        RECT 2.904000 0.395000 2.965000 0.727000 ;
        RECT 2.719000 0.267000 2.780000 0.435000 ;
        RECT 2.596000 0.390000 2.657000 0.852000 ;
        RECT 2.287000 0.163000 2.348000 0.445000 ;
        RECT 1.803000 0.614000 1.864000 0.701000 ;
        RECT 1.611000 0.424000 1.672000 0.564000 ;
        RECT 1.415000 0.249000 1.476000 0.701000 ;
        RECT 1.388000 0.646000 1.449000 0.792000 ;
        RECT 1.135000 0.856000 1.196000 0.962000 ;
        RECT 0.675000 0.856000 0.736000 0.993000 ;
        RECT 0.552000 0.732000 0.613000 0.860000 ;
        RECT 0.044000 0.317000 0.105000 0.769000 ;
        RECT 2.857000 0.206000 3.141000 0.263000 ;
        RECT 3.779000 0.407000 4.184000 0.462000 ;
        RECT 3.497000 0.583000 4.088000 0.638000 ;
        RECT 3.299000 0.362000 3.479000 0.417000 ;
        RECT 2.925000 0.802000 3.141000 0.857000 ;
        RECT 2.857000 0.206000 3.840000 0.261000 ;
        RECT 2.719000 0.380000 2.843000 0.435000 ;
        RECT 2.287000 0.390000 2.657000 0.445000 ;
        RECT 2.185000 0.939000 3.559000 0.994000 ;
        RECT 2.123000 0.501000 2.535000 0.556000 ;
        RECT 1.987000 0.501000 2.473000 0.556000 ;
        RECT 1.925000 0.501000 2.472000 0.556000 ;
        RECT 1.856000 0.163000 2.348000 0.218000 ;
        RECT 1.611000 0.424000 1.987000 0.479000 ;
        RECT 1.388000 0.646000 1.864000 0.701000 ;
        RECT 1.323000 0.249000 1.476000 0.304000 ;
        RECT 1.257000 0.890000 1.549000 0.945000 ;
        RECT 0.675000 0.856000 1.196000 0.911000 ;
        RECT 0.552000 0.732000 1.319000 0.787000 ;
        RECT 0.533000 0.938000 0.736000 0.993000 ;
        RECT 0.429000 0.608000 0.691000 0.663000 ;
        RECT 0.384000 0.206000 1.200000 0.261000 ;
        RECT 0.077000 0.805000 0.613000 0.860000 ;
        RECT 2.629000 0.267000 2.780000 0.321000 ;
        RECT 2.381000 0.798000 2.657000 0.852000 ;
        RECT 0.557000 0.348000 0.911000 0.402000 ;
        RECT 0.557000 0.348000 0.912000 0.398000 ;
        RECT 0.600000 0.348000 0.649000 0.676000 ;
        RECT 2.927000 0.382000 2.965000 0.727000 ;
        RECT 1.415000 0.249000 1.449000 0.792000 ;
        RECT 3.527000 0.526000 3.559000 1.020000 ;
        RECT 2.185000 0.614000 2.213000 0.994000 ;
        RECT 0.077000 0.317000 0.105000 0.860000 ;
        RECT 1.925000 0.398000 1.949000 0.876000 ;
        RECT 2.719000 0.240000 2.720000 0.435000 ;
    END
END SDFFRHQX1

MACRO OAI221XL
    CLASS CORE ;
    FOREIGN OAI221XL 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.300000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.336000 0.642000 0.519000 0.779000 ;
        RECT 0.421000 0.640000 0.516000 0.779000 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.622000 0.639000 0.718000 0.755000 ;
        RECT 0.803000 0.700000 0.868000 0.761000 ;
        RECT 0.622000 0.700000 0.868000 0.755000 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.187000 0.433000 0.359000 0.550000 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.039000 0.640000 0.146000 0.821000 ;
        END
    END B1
    PIN C0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.968000 0.521000 1.075000 0.654000 ;
        END
    END C0
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.300000 1.280000 ;
        RECT 0.681000 1.078000 0.777000 1.280000 ;
        RECT 0.051000 1.078000 0.146000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.300000 0.080000 ;
        RECT 0.366000 -0.080000 0.461000 0.122000 ;
        RECT 0.051000 -0.080000 0.146000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.095000 0.258000 1.240000 0.339000 ;
        RECT 0.895000 0.865000 0.990000 0.946000 ;
        RECT 0.366000 0.865000 0.461000 0.946000 ;
        RECT 1.175000 0.258000 1.240000 0.920000 ;
        RECT 0.366000 0.865000 1.240000 0.920000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.722000 0.339000 0.817000 0.420000 ;
        RECT 0.208000 0.252000 0.304000 0.333000 ;
        RECT 0.722000 0.252000 0.786000 0.420000 ;
        RECT 0.208000 0.252000 0.786000 0.307000 ;
    END
END OAI221XL

MACRO OAI21XL
    CLASS CORE ;
    FOREIGN OAI21XL 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 0.700000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.212000 0.479000 0.388000 0.571000 ;
        RECT 0.232000 0.439000 0.293000 0.571000 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.048000 0.433000 0.138000 0.618000 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.387000 0.640000 0.528000 0.767000 ;
        END
    END B0
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 0.700000 1.280000 ;
        RECT 0.536000 1.078000 0.626000 1.280000 ;
        RECT 0.048000 0.910000 0.138000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 0.700000 0.080000 ;
        RECT 0.196000 -0.080000 0.286000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.387000 0.848000 0.477000 0.929000 ;
        RECT 0.589000 0.439000 0.650000 0.915000 ;
        RECT 0.582000 0.161000 0.643000 0.494000 ;
        RECT 0.582000 0.439000 0.650000 0.494000 ;
        RECT 0.589000 0.161000 0.643000 0.915000 ;
        RECT 0.546000 0.161000 0.643000 0.215000 ;
        RECT 0.387000 0.861000 0.650000 0.915000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.398000 0.332000 0.488000 0.413000 ;
        RECT 0.048000 0.296000 0.138000 0.377000 ;
        RECT 0.398000 0.296000 0.459000 0.413000 ;
        RECT 0.048000 0.296000 0.459000 0.351000 ;
    END
END OAI21XL

MACRO NOR4BX1
    CLASS CORE ;
    FOREIGN NOR4BX1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.100000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN AN
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.038000 0.395000 0.144000 0.531000 ;
        RECT 0.049000 0.395000 0.143000 0.532000 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.697000 0.413000 0.878000 0.513000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.508000 0.557000 0.603000 0.638000 ;
        RECT 0.464000 0.439000 0.528000 0.612000 ;
        RECT 0.464000 0.557000 0.603000 0.612000 ;
        RECT 0.426000 0.439000 0.528000 0.494000 ;
        RECT 0.508000 0.439000 0.528000 0.638000 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.336000 0.556000 0.400000 0.755000 ;
        RECT 0.243000 0.700000 0.307000 0.761000 ;
        RECT 0.243000 0.700000 0.400000 0.755000 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.100000 1.280000 ;
        RECT 0.233000 1.078000 0.328000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.100000 0.080000 ;
        RECT 0.583000 -0.080000 0.678000 0.122000 ;
        RECT 0.233000 -0.080000 0.328000 0.122000 ;
        RECT 0.950000 -0.080000 1.044000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.917000 0.718000 1.036000 0.799000 ;
        RECT 0.428000 0.262000 0.889000 0.343000 ;
        RECT 0.972000 0.288000 1.036000 0.799000 ;
        RECT 0.972000 0.439000 1.040000 0.494000 ;
        RECT 0.428000 0.288000 1.036000 0.343000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.050000 0.707000 0.144000 0.788000 ;
        RECT 0.050000 0.246000 0.144000 0.327000 ;
        RECT 0.667000 0.594000 0.731000 0.876000 ;
        RECT 0.208000 0.273000 0.272000 0.643000 ;
        RECT 0.081000 0.588000 0.144000 0.876000 ;
        RECT 0.667000 0.594000 0.908000 0.649000 ;
        RECT 0.081000 0.821000 0.731000 0.876000 ;
        RECT 0.081000 0.588000 0.272000 0.643000 ;
        RECT 0.050000 0.273000 0.272000 0.327000 ;
    END
END NOR4BX1

MACRO NOR3X1
    CLASS CORE ;
    FOREIGN NOR3X1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 0.700000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.456000 0.536000 0.546000 0.617000 ;
        RECT 0.456000 0.536000 0.517000 0.761000 ;
        RECT 0.407000 0.706000 0.517000 0.761000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.232000 0.421000 0.361000 0.561000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.048000 0.536000 0.137000 0.694000 ;
        RECT 0.048000 0.536000 0.138000 0.617000 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 0.700000 1.280000 ;
        RECT 0.048000 0.900000 0.138000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 0.700000 0.080000 ;
        RECT 0.345000 -0.080000 0.435000 0.122000 ;
        RECT 0.048000 -0.080000 0.138000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.557000 0.839000 0.666000 0.924000 ;
        RECT 0.196000 0.269000 0.668000 0.350000 ;
        RECT 0.607000 0.269000 0.668000 0.894000 ;
        RECT 0.607000 0.269000 0.666000 0.924000 ;
        RECT 0.557000 0.839000 0.668000 0.894000 ;
        END
    END Y
END NOR3X1

MACRO NOR2BX1
    CLASS CORE ;
    FOREIGN NOR2BX1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 0.700000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN AN
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.037000 0.486000 0.138000 0.633000 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.321000 0.567000 0.411000 0.670000 ;
        RECT 0.321000 0.567000 0.525000 0.633000 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 0.700000 1.280000 ;
        RECT 0.212000 0.916000 0.302000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 0.700000 0.080000 ;
        RECT 0.562000 -0.080000 0.652000 0.122000 ;
        RECT 0.263000 -0.080000 0.353000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.562000 0.706000 0.666000 0.858000 ;
        RECT 0.411000 0.269000 0.501000 0.350000 ;
        RECT 0.605000 0.295000 0.666000 0.858000 ;
        RECT 0.411000 0.295000 0.666000 0.350000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.461000 0.430000 0.544000 0.511000 ;
        RECT 0.048000 0.715000 0.138000 0.796000 ;
        RECT 0.048000 0.304000 0.138000 0.385000 ;
        RECT 0.048000 0.323000 0.260000 0.385000 ;
        RECT 0.199000 0.323000 0.260000 0.770000 ;
        RECT 0.260000 0.443000 0.461000 0.498000 ;
        RECT 0.048000 0.715000 0.260000 0.770000 ;
    END
END NOR2BX1

MACRO NOR2X1
    CLASS CORE ;
    FOREIGN NOR2X1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 0.600000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.242000 0.407000 0.421000 0.502000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.061000 0.548000 0.164000 0.643000 ;
        RECT 0.042000 0.567000 0.255000 0.643000 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 0.600000 1.280000 ;
        RECT 0.055000 1.078000 0.158000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 0.600000 0.080000 ;
        RECT 0.442000 -0.080000 0.545000 0.122000 ;
        RECT 0.055000 -0.080000 0.158000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.442000 0.626000 0.561000 0.774000 ;
        RECT 0.248000 0.269000 0.352000 0.350000 ;
        RECT 0.491000 0.295000 0.561000 0.774000 ;
        RECT 0.248000 0.295000 0.561000 0.350000 ;
        END
    END Y
END NOR2X1

MACRO NAND4BBX1
    CLASS CORE ;
    FOREIGN NAND4BBX1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.400000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN AN
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.070000 0.498000 1.188000 0.633000 ;
        RECT 1.070000 0.498000 1.201000 0.579000 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.041000 0.433000 0.142000 0.574000 ;
        END
    END BN
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.502000 0.555000 0.610000 0.636000 ;
        RECT 0.549000 0.439000 0.610000 0.636000 ;
        RECT 0.549000 0.439000 0.643000 0.494000 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.327000 0.519000 0.412000 0.600000 ;
        RECT 0.351000 0.439000 0.412000 0.600000 ;
        RECT 0.351000 0.439000 0.468000 0.494000 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.400000 1.280000 ;
        RECT 0.957000 1.078000 1.077000 1.280000 ;
        RECT 0.607000 1.078000 0.697000 1.280000 ;
        RECT 0.247000 1.078000 0.337000 1.280000 ;
        RECT 0.261000 1.065000 0.322000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.098000 -0.080000 0.316000 0.122000 ;
        RECT 0.000000 -0.080000 1.400000 0.080000 ;
        RECT 1.262000 -0.080000 1.352000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.788000 0.742000 0.878000 0.839000 ;
        RECT 0.737000 0.755000 0.878000 0.839000 ;
        RECT 1.262000 0.201000 1.343000 0.306000 ;
        RECT 0.874000 0.201000 0.964000 0.282000 ;
        RECT 0.427000 0.742000 0.517000 0.823000 ;
        RECT 0.427000 0.742000 0.582000 0.810000 ;
        RECT 1.306000 0.573000 1.367000 0.933000 ;
        RECT 1.282000 0.201000 1.343000 0.627000 ;
        RECT 0.817000 0.742000 0.878000 0.933000 ;
        RECT 0.874000 0.201000 1.343000 0.256000 ;
        RECT 0.427000 0.755000 0.878000 0.810000 ;
        RECT 1.282000 0.573000 1.367000 0.627000 ;
        RECT 0.817000 0.879000 1.367000 0.933000 ;
        RECT 1.306000 0.201000 1.343000 0.933000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 1.059000 0.311000 1.149000 0.392000 ;
        RECT 0.890000 0.419000 1.005000 0.500000 ;
        RECT 0.709000 0.555000 0.799000 0.636000 ;
        RECT 0.048000 0.746000 0.138000 0.827000 ;
        RECT 0.048000 0.293000 0.138000 0.374000 ;
        RECT 0.944000 0.337000 1.005000 0.810000 ;
        RECT 0.738000 0.302000 0.799000 0.636000 ;
        RECT 0.203000 0.302000 0.264000 0.801000 ;
        RECT 0.944000 0.755000 1.245000 0.810000 ;
        RECT 0.944000 0.337000 1.149000 0.392000 ;
        RECT 0.203000 0.302000 0.799000 0.357000 ;
        RECT 0.048000 0.746000 0.264000 0.801000 ;
        RECT 0.048000 0.302000 0.709000 0.357000 ;
    END
END NAND4BBX1

MACRO NAND3BX2
    CLASS CORE ;
    FOREIGN NAND3BX2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.400000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN AN
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.262000 0.467000 1.363000 0.594000 ;
        RECT 1.267000 0.433000 1.358000 0.594000 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.737000 0.433000 0.838000 0.604000 ;
        RECT 0.355000 0.514000 0.445000 0.604000 ;
        RECT 0.737000 0.507000 0.870000 0.588000 ;
        RECT 0.355000 0.549000 0.838000 0.604000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.082000 0.439000 0.172000 0.573000 ;
        RECT 0.957000 0.462000 1.047000 0.543000 ;
        RECT 0.972000 0.462000 1.033000 0.881000 ;
        RECT 0.111000 0.439000 0.172000 0.881000 ;
        RECT 0.111000 0.826000 1.033000 0.881000 ;
        RECT 0.057000 0.439000 0.172000 0.494000 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.400000 1.280000 ;
        RECT 1.058000 0.952000 1.148000 1.280000 ;
        RECT 0.471000 0.952000 0.561000 1.280000 ;
        RECT 0.102000 0.952000 0.192000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.400000 0.080000 ;
        RECT 1.055000 -0.080000 1.161000 0.122000 ;
        RECT 1.055000 -0.080000 1.145000 0.247000 ;
        RECT 0.064000 -0.080000 0.154000 0.247000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.651000 0.689000 0.741000 0.770000 ;
        RECT 0.567000 0.164000 0.658000 0.245000 ;
        RECT 0.282000 0.689000 0.373000 0.770000 ;
        RECT 0.643000 0.689000 0.741000 0.767000 ;
        RECT 0.233000 0.689000 0.407000 0.767000 ;
        RECT 0.233000 0.700000 0.741000 0.767000 ;
        RECT 0.233000 0.177000 0.294000 0.767000 ;
        RECT 0.233000 0.177000 0.658000 0.232000 ;
        RECT 0.282000 0.177000 0.294000 0.770000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 1.262000 0.279000 1.352000 0.379000 ;
        RECT 1.262000 0.702000 1.352000 0.783000 ;
        RECT 0.567000 0.410000 0.658000 0.490000 ;
        RECT 1.140000 0.324000 1.201000 0.757000 ;
        RECT 0.597000 0.324000 0.658000 0.490000 ;
        RECT 1.140000 0.702000 1.352000 0.757000 ;
        RECT 0.597000 0.324000 1.352000 0.379000 ;
    END
END NAND3BX2

MACRO NAND3X1
    CLASS CORE ;
    FOREIGN NAND3X1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 0.700000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.439000 0.501000 0.529000 0.582000 ;
        RECT 0.439000 0.306000 0.500000 0.582000 ;
        RECT 0.407000 0.306000 0.500000 0.361000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.232000 0.544000 0.349000 0.676000 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.050000 0.425000 0.141000 0.590000 ;
        END
    END C
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.048000 1.078000 0.483000 1.280000 ;
        RECT 0.000000 1.120000 0.700000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 0.700000 0.080000 ;
        RECT 0.064000 -0.080000 0.154000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.562000 0.167000 0.652000 0.307000 ;
        RECT 0.562000 0.731000 0.655000 0.812000 ;
        RECT 0.203000 0.731000 0.293000 0.812000 ;
        RECT 0.581000 0.695000 0.655000 0.812000 ;
        RECT 0.591000 0.167000 0.652000 0.812000 ;
        RECT 0.203000 0.744000 0.655000 0.799000 ;
        END
    END Y
END NAND3X1

MACRO NAND2BX1
    CLASS CORE ;
    FOREIGN NAND2BX1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 0.700000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN AN
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.056000 0.901000 0.196000 1.033000 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.232000 0.439000 0.377000 0.545000 ;
        RECT 0.212000 0.461000 0.391000 0.545000 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.377000 1.078000 0.636000 1.280000 ;
        RECT 0.000000 1.120000 0.700000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 0.700000 0.080000 ;
        RECT 0.207000 -0.080000 0.297000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.557000 0.289000 0.647000 0.370000 ;
        RECT 0.467000 0.300000 0.647000 0.367000 ;
        RECT 0.586000 0.289000 0.647000 0.808000 ;
        RECT 0.407000 0.306000 0.647000 0.361000 ;
        RECT 0.398000 0.754000 0.647000 0.808000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.048000 0.740000 0.138000 0.821000 ;
        RECT 0.048000 0.274000 0.138000 0.355000 ;
        RECT 0.463000 0.605000 0.524000 0.694000 ;
        RECT 0.062000 0.274000 0.123000 0.821000 ;
        RECT 0.138000 0.605000 0.524000 0.660000 ;
        RECT 0.123000 0.605000 0.463000 0.660000 ;
        RECT 0.062000 0.605000 0.138000 0.660000 ;
    END
END NAND2BX1

MACRO NAND2X1
    CLASS CORE ;
    FOREIGN NAND2X1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 0.600000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.242000 0.530000 0.421000 0.633000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.042000 0.438000 0.158000 0.598000 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.055000 1.078000 0.359000 1.280000 ;
        RECT 0.000000 1.120000 0.600000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 0.600000 0.080000 ;
        RECT 0.055000 -0.080000 0.158000 0.328000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.442000 0.282000 0.545000 0.367000 ;
        RECT 0.248000 0.688000 0.352000 0.769000 ;
        RECT 0.494000 0.300000 0.564000 0.743000 ;
        RECT 0.442000 0.300000 0.564000 0.367000 ;
        RECT 0.248000 0.688000 0.564000 0.743000 ;
        RECT 0.494000 0.282000 0.545000 0.743000 ;
        END
    END Y
END NAND2X1

MACRO MXI2X1
    CLASS CORE ;
    FOREIGN MXI2X1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.300000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.128000 0.433000 1.261000 0.543000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.411000 0.433000 0.529000 0.555000 ;
        END
    END B
    PIN S0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.198000 0.524000 0.332000 0.633000 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.300000 1.280000 ;
        RECT 1.152000 1.064000 1.251000 1.280000 ;
        RECT 0.304000 0.954000 0.400000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.300000 0.080000 ;
        RECT 1.151000 -0.080000 1.247000 0.122000 ;
        RECT 0.315000 -0.080000 0.411000 0.347000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.764000 0.573000 0.868000 0.805000 ;
        RECT 0.748000 0.724000 0.868000 0.805000 ;
        RECT 0.748000 0.281000 0.844000 0.362000 ;
        RECT 0.764000 0.281000 0.829000 0.805000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.049000 0.736000 0.152000 0.870000 ;
        RECT 0.049000 0.292000 0.163000 0.381000 ;
        RECT 0.962000 0.279000 1.058000 0.360000 ;
        RECT 0.590000 0.933000 0.698000 1.014000 ;
        RECT 0.535000 0.281000 0.677000 0.362000 ;
        RECT 0.529000 0.679000 0.677000 0.760000 ;
        RECT 0.974000 0.710000 1.069000 0.790000 ;
        RECT 0.049000 0.292000 0.165000 0.368000 ;
        RECT 0.975000 0.279000 1.040000 0.790000 ;
        RECT 0.612000 0.281000 0.677000 0.760000 ;
        RECT 0.049000 0.292000 0.114000 0.870000 ;
        RECT 0.590000 0.815000 0.654000 1.014000 ;
        RECT 0.049000 0.815000 0.654000 0.870000 ;
    END
END MXI2X1

MACRO MX2X1
    CLASS CORE ;
    FOREIGN MX2X1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.400000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.000000 0.433000 1.188000 0.527000 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.292000 0.635000 0.387000 0.767000 ;
        RECT 0.292000 0.688000 0.488000 0.767000 ;
        END
    END B
    PIN S0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.037000 0.944000 0.188000 1.033000 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.400000 1.280000 ;
        RECT 1.050000 1.078000 1.140000 1.280000 ;
        RECT 0.249000 0.852000 0.339000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.400000 0.080000 ;
        RECT 1.049000 -0.080000 1.139000 0.122000 ;
        RECT 0.264000 -0.080000 0.349000 0.342000 ;
        RECT 0.261000 0.291000 0.351000 0.342000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.198000 0.754000 1.363000 0.946000 ;
        RECT 1.250000 0.268000 1.363000 0.379000 ;
        RECT 1.248000 0.268000 1.363000 0.361000 ;
        RECT 1.302000 0.268000 1.363000 0.946000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.671000 0.789000 0.793000 0.882000 ;
        RECT 0.460000 0.508000 0.546000 0.599000 ;
        RECT 1.103000 0.615000 1.193000 0.696000 ;
        RECT 0.463000 0.269000 0.553000 0.350000 ;
        RECT 0.048000 0.752000 0.138000 0.833000 ;
        RECT 0.048000 0.276000 0.138000 0.357000 ;
        RECT 1.035000 0.621000 1.193000 0.696000 ;
        RECT 1.035000 0.621000 1.096000 0.968000 ;
        RECT 0.862000 0.269000 0.923000 0.838000 ;
        RECT 0.732000 0.280000 0.793000 0.968000 ;
        RECT 0.610000 0.393000 0.671000 0.720000 ;
        RECT 0.549000 0.665000 0.610000 0.887000 ;
        RECT 0.492000 0.269000 0.553000 0.448000 ;
        RECT 0.062000 0.276000 0.123000 0.833000 ;
        RECT 0.732000 0.913000 1.096000 0.968000 ;
        RECT 0.654000 0.280000 0.793000 0.335000 ;
        RECT 0.549000 0.665000 0.671000 0.720000 ;
        RECT 0.492000 0.393000 0.671000 0.448000 ;
        RECT 0.440000 0.832000 0.610000 0.887000 ;
        RECT 0.138000 0.524000 0.546000 0.579000 ;
        RECT 0.123000 0.524000 0.460000 0.579000 ;
        RECT 0.062000 0.524000 0.440000 0.579000 ;
    END
END MX2X1

MACRO INVXL
    CLASS CORE ;
    FOREIGN INVXL 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 0.400000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.042000 0.433000 0.158000 0.598000 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 0.400000 1.280000 ;
        RECT 0.155000 0.925000 0.258000 1.280000 ;
        RECT 0.083000 0.925000 0.329000 0.975000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.055000 -0.080000 0.300000 0.122000 ;
        RECT 0.000000 -0.080000 0.400000 0.080000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.242000 0.567000 0.358000 0.768000 ;
        RECT 0.236000 0.321000 0.339000 0.439000 ;
        RECT 0.242000 0.321000 0.312000 0.768000 ;
        END
    END Y
END INVXL

MACRO INVX2
    CLASS CORE ;
    FOREIGN INVX2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 0.600000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.150000 0.433000 0.395000 0.574000 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 0.600000 1.280000 ;
        RECT 0.394000 1.078000 0.497000 1.280000 ;
        RECT 0.395000 1.064000 0.495000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 0.600000 0.080000 ;
        RECT 0.164000 -0.080000 0.267000 0.361000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.442000 0.183000 0.558000 0.376000 ;
        RECT 0.224000 0.661000 0.327000 0.854000 ;
        RECT 0.465000 0.627000 0.558000 0.715000 ;
        RECT 0.488000 0.183000 0.558000 0.715000 ;
        RECT 0.224000 0.661000 0.558000 0.715000 ;
        END
    END Y
END INVX2

MACRO INVX1
    CLASS CORE ;
    FOREIGN INVX1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 0.400000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.042000 0.433000 0.173000 0.568000 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 0.400000 1.280000 ;
        RECT 0.055000 1.078000 0.158000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 0.400000 0.080000 ;
        RECT 0.055000 -0.080000 0.158000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.242000 0.564000 0.358000 0.848000 ;
        RECT 0.253000 0.321000 0.323000 0.848000 ;
        END
    END Y
END INVX1

MACRO BUFX2
    CLASS CORE ;
    FOREIGN BUFX2 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 0.700000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.037000 0.418000 0.236000 0.538000 ;
        END
    END A
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 0.700000 1.280000 ;
        RECT 0.223000 1.078000 0.313000 1.280000 ;
        RECT 0.237000 1.065000 0.298000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 0.700000 0.080000 ;
        RECT 0.233000 -0.080000 0.323000 0.122000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.435000 0.331000 0.525000 0.412000 ;
        RECT 0.424000 0.655000 0.514000 0.736000 ;
        RECT 0.562000 0.357000 0.623000 0.710000 ;
        RECT 0.562000 0.439000 0.643000 0.494000 ;
        RECT 0.435000 0.357000 0.623000 0.412000 ;
        RECT 0.424000 0.655000 0.623000 0.710000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.302000 0.490000 0.430000 0.571000 ;
        RECT 0.074000 0.657000 0.164000 0.738000 ;
        RECT 0.074000 0.275000 0.164000 0.356000 ;
        RECT 0.302000 0.301000 0.363000 0.712000 ;
        RECT 0.074000 0.657000 0.363000 0.712000 ;
        RECT 0.074000 0.301000 0.363000 0.356000 ;
    END
END BUFX2

MACRO AOI32X1
    CLASS CORE ;
    FOREIGN AOI32X1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.300000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.411000 0.383000 0.597000 0.500000 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.246000 0.571000 0.416000 0.680000 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.039000 0.400000 0.225000 0.500000 ;
        END
    END A2
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.712000 0.560000 0.889000 0.640000 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.877000 0.381000 1.054000 0.494000 ;
        END
    END B1
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 1.300000 1.280000 ;
        RECT 0.456000 0.925000 0.552000 1.280000 ;
        RECT 0.051000 0.800000 0.146000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 1.300000 0.080000 ;
        RECT 0.948000 -0.080000 1.044000 0.122000 ;
        RECT 0.066000 -0.080000 0.131000 0.325000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.154000 0.223000 1.240000 0.306000 ;
        RECT 1.175000 0.223000 1.240000 0.820000 ;
        RECT 0.861000 0.765000 1.240000 0.820000 ;
        RECT 0.568000 0.223000 1.240000 0.277000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.674000 0.800000 0.739000 0.963000 ;
        RECT 0.674000 0.908000 1.159000 0.963000 ;
        RECT 0.253000 0.800000 0.739000 0.855000 ;
    END
END AOI32X1

MACRO AOI22X1
    CLASS CORE ;
    FOREIGN AOI22X1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 0.900000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.499000 0.394000 0.592000 0.475000 ;
        RECT 0.419000 0.407000 0.592000 0.475000 ;
        RECT 0.419000 0.407000 0.481000 0.494000 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.577000 0.538000 0.731000 0.633000 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.239000 0.567000 0.415000 0.663000 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.052000 0.421000 0.145000 0.589000 ;
        END
    END B1
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 0.900000 1.280000 ;
        RECT 0.229000 1.078000 0.322000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 0.900000 0.080000 ;
        RECT 0.758000 -0.080000 0.851000 0.122000 ;
        RECT 0.049000 -0.080000 0.142000 0.330000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.779000 0.265000 0.862000 0.361000 ;
        RECT 0.584000 0.699000 0.676000 0.780000 ;
        RECT 0.398000 0.252000 0.491000 0.333000 ;
        RECT 0.799000 0.265000 0.862000 0.754000 ;
        RECT 0.584000 0.699000 0.862000 0.754000 ;
        RECT 0.398000 0.265000 0.862000 0.320000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.049000 0.726000 0.142000 0.933000 ;
        RECT 0.758000 0.854000 0.851000 0.935000 ;
        RECT 0.409000 0.865000 0.502000 0.946000 ;
        RECT 0.409000 0.880000 0.851000 0.935000 ;
        RECT 0.049000 0.879000 0.502000 0.933000 ;
        RECT 0.049000 0.880000 0.851000 0.933000 ;
    END
END AOI22X1

MACRO AOI21X1
    CLASS CORE ;
    FOREIGN AOI21X1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 0.700000 BY 1.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ; 
    PIN A0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.232000 0.306000 0.293000 0.623000 ;
        RECT 0.232000 0.568000 0.379000 0.623000 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.050000 0.492000 0.141000 0.615000 ;
        RECT 0.050000 0.433000 0.138000 0.615000 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.477000 0.439000 0.542000 0.627000 ;
        RECT 0.407000 0.439000 0.542000 0.494000 ;
        END
    END B0
    PIN VDD
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE POWER ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 1.120000 0.700000 1.280000 ;
        RECT 0.217000 0.852000 0.308000 1.280000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        SHAPE ABUTMENT ;
        USE GROUND ;
        PORT
        LAYER Metal1 ;
        RECT 0.000000 -0.080000 0.700000 0.080000 ;
        RECT 0.536000 -0.080000 0.626000 0.122000 ;
        RECT 0.048000 -0.080000 0.138000 0.334000 ;
        END
    END VSS
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 0.582000 0.706000 0.664000 0.940000 ;
        RECT 0.387000 0.295000 0.477000 0.376000 ;
        RECT 0.557000 0.860000 0.664000 0.940000 ;
        RECT 0.603000 0.321000 0.664000 0.940000 ;
        RECT 0.387000 0.321000 0.664000 0.376000 ;
        END
    END Y
    OBS
        LAYER Metal1 ;
        RECT 0.048000 0.696000 0.477000 0.751000 ;
    END
END AOI21X1

MACRO PDIDGZ
    CLASS PAD ;
    FOREIGN PDIDGZ 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 4.000000 BY 23.500000 ;
    SYMMETRY X Y R90 ;
    SITE CoreSite ; 
    PIN C
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 3.217000 23.400000 3.417000 23.500000 ;
        LAYER Metal2 ;
        RECT 3.217000 23.400000 3.417000 23.500000 ;
        LAYER Metal3 ;
        RECT 3.217000 23.400000 3.417000 23.500000 ;
        LAYER Metal4 ;
        RECT 3.217000 23.400000 3.417000 23.500000 ;
        LAYER Metal5 ;
        RECT 3.217000 23.400000 3.417000 23.500000 ;
        END
    END C
    PIN PAD
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.877000 0.000000 2.224000 0.136000 ;
        LAYER Metal2 ;
        RECT 1.877000 0.000000 2.224000 0.136000 ;
        END
    END PAD
    OBS
        LAYER Metal1 ;
        RECT 0.000000 0.196000 3.167000 23.500000 ;
        RECT 0.000000 0.000000 1.827000 23.500000 ;
        RECT 2.274000 0.000000 4.000000 23.350000 ;
        RECT 2.274000 0.000000 3.167000 23.500000 ;
        RECT 3.467000 0.000000 4.000000 23.500000 ;
        LAYER Via1 ;
        RECT 0.000000 0.000000 4.000000 23.500000 ;
        LAYER Metal2 ;
        RECT 0.000000 0.196000 3.167000 23.500000 ;
        RECT 0.000000 0.000000 1.827000 23.500000 ;
        RECT 2.274000 0.000000 4.000000 23.350000 ;
        RECT 2.274000 0.000000 3.167000 23.500000 ;
        RECT 3.467000 0.000000 4.000000 23.500000 ;
        LAYER Via2 ;
        RECT 0.000000 0.000000 4.000000 23.500000 ;
        LAYER Metal3 ;
        RECT 0.000000 0.000000 4.000000 23.350000 ;
        RECT 0.000000 0.000000 3.167000 23.500000 ;
        RECT 3.467000 0.000000 4.000000 23.500000 ;
        LAYER Via3 ;
        RECT 0.000000 0.000000 4.000000 23.500000 ;
        LAYER Metal4 ;
        RECT 0.000000 0.000000 4.000000 23.350000 ;
        RECT 0.000000 0.000000 3.167000 23.500000 ;
        RECT 3.467000 0.000000 4.000000 23.500000 ;
        LAYER Via4 ;
        RECT 0.000000 0.000000 4.000000 23.500000 ;
        LAYER Metal5 ;
        RECT 0.000000 0.000000 4.000000 23.350000 ;
        RECT 0.000000 0.000000 3.167000 23.500000 ;
        RECT 3.467000 0.000000 4.000000 23.500000 ;
        LAYER Via5 ;
        RECT 0.000000 0.000000 4.000000 23.500000 ;
        LAYER Metal6 ;
        RECT 0.000000 0.000000 4.000000 23.500000 ;
    END
END PDIDGZ

MACRO PDO04CDG
    CLASS PAD ;
    FOREIGN PDO04CDG 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 4.000000 BY 23.500000 ;
    SYMMETRY X Y R90 ;
    SITE CoreSite ; 
    PIN I
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 3.217000 23.400000 3.417000 23.500000 ;
        LAYER Metal2 ;
        RECT 3.217000 23.400000 3.417000 23.500000 ;
        LAYER Metal3 ;
        RECT 3.217000 23.400000 3.417000 23.500000 ;
        LAYER Metal4 ;
        RECT 3.217000 23.400000 3.417000 23.500000 ;
        LAYER Metal5 ;
        RECT 3.217000 23.400000 3.417000 23.500000 ;
        END
    END I
    PIN PAD
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER Metal1 ;
        RECT 1.877000 0.000000 2.224000 0.136000 ;
        LAYER Metal2 ;
        RECT 1.877000 0.000000 2.224000 0.136000 ;
        END
    END PAD
    OBS
        LAYER Metal1 ;
        RECT 0.000000 0.196000 3.167000 23.500000 ;
        RECT 0.000000 0.000000 1.827000 23.500000 ;
        RECT 2.274000 0.000000 4.000000 23.350000 ;
        RECT 2.274000 0.000000 3.167000 23.500000 ;
        RECT 3.467000 0.000000 4.000000 23.500000 ;
        LAYER Via1 ;
        RECT 0.000000 0.000000 4.000000 23.500000 ;
        LAYER Metal2 ;
        RECT 0.000000 0.196000 3.167000 23.500000 ;
        RECT 0.000000 0.000000 1.827000 23.500000 ;
        RECT 2.274000 0.000000 4.000000 23.350000 ;
        RECT 2.274000 0.000000 3.167000 23.500000 ;
        RECT 3.467000 0.000000 4.000000 23.500000 ;
        LAYER Via2 ;
        RECT 0.000000 0.000000 4.000000 23.500000 ;
        LAYER Metal3 ;
        RECT 0.000000 0.000000 4.000000 23.350000 ;
        RECT 0.000000 0.000000 3.167000 23.500000 ;
        RECT 3.467000 0.000000 4.000000 23.500000 ;
        LAYER Via3 ;
        RECT 0.000000 0.000000 4.000000 23.500000 ;
        LAYER Metal4 ;
        RECT 0.000000 0.000000 4.000000 23.350000 ;
        RECT 0.000000 0.000000 3.167000 23.500000 ;
        RECT 3.467000 0.000000 4.000000 23.500000 ;
        LAYER Via4 ;
        RECT 0.000000 0.000000 4.000000 23.500000 ;
        LAYER Metal5 ;
        RECT 0.000000 0.000000 4.000000 23.350000 ;
        RECT 0.000000 0.000000 3.167000 23.500000 ;
        RECT 3.467000 0.000000 4.000000 23.500000 ;
        LAYER Via5 ;
        RECT 0.000000 0.000000 4.000000 23.500000 ;
        LAYER Metal6 ;
        RECT 0.000000 0.000000 4.000000 23.500000 ;
    END
END PDO04CDG

END LIBRARY

