VERSION 5.7 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS	2000 ;
END UNITS

MANUFACTURINGGRID	0.0025 ;

SITE core
  SIZE 0.19 BY 1.71 ;
  CLASS CORE ;
END core

LAYER metal1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.19 ;
  WIDTH 0.065 ;
END metal1

LAYER metal2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.19 ;
  WIDTH 0.07 ;
END metal2

LAYER metal3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.19 ;
  WIDTH 0.07 ;
END metal3

LAYER metal4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.285 ;
  WIDTH 0.14 ;
END metal4

MACRO INV_X1
    CLASS CORE ;
    FOREIGN INV_X1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.760 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.465 0.150 0.53 1.255 ;
        RECT 0.415 0.150 0.61 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.210 0.340 0.34 0.405 ;
        END
    END a
END INV_X1

MACRO INV_X2
    CLASS CORE ;
    FOREIGN INV_X2 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.520 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.925 0.150 1.12 1.255 ;
        RECT 0.835 0.150 1.225 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.420 0.340 0.68 0.405 ;
        END
    END a
END INV_X2

MACRO INV_X3
    CLASS CORE ;
    FOREIGN INV_X3 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.900 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.160 0.150 1.355 1.255 ;
        RECT 1.040 0.150 1.495 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.525 0.340 0.85 0.405 ;
        END
    END a
END INV_X3

MACRO INV_X4
    CLASS CORE ;
    FOREIGN INV_X4 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.900 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.160 0.150 1.355 1.255 ;
        RECT 1.040 0.150 1.495 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.525 0.340 0.85 0.405 ;
        END
    END a
END INV_X4

MACRO INV_X6
    CLASS CORE ;
    FOREIGN INV_X6 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.280 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.150 1.65 1.255 ;
        RECT 1.250 0.150 1.77 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.630 0.340 1.02 0.405 ;
        END
    END a
END INV_X6

MACRO INV_X8
    CLASS CORE ;
    FOREIGN INV_X8 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.620 0.150 1.945 1.255 ;
        RECT 1.460 0.150 2.11 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.735 0.340 1.19 0.405 ;
        END
    END a
END INV_X8

MACRO INV_X10
    CLASS CORE ;
    FOREIGN INV_X10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.620 0.150 1.945 1.255 ;
        RECT 1.460 0.150 2.11 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.735 0.340 1.19 0.405 ;
        END
    END a
END INV_X10

MACRO INV_X20
    CLASS CORE ;
    FOREIGN INV_X20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.315 0.150 2.77 1.255 ;
        RECT 2.085 0.150 2.995 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.050 0.340 1.7 0.405 ;
        END
    END a
END INV_X20

MACRO INV_X40
    CLASS CORE ;
    FOREIGN INV_X40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.940 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.010 0.150 3.595 1.255 ;
        RECT 2.710 0.150 3.88 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.365 0.340 2.21 0.405 ;
        END
    END a
END INV_X40

MACRO INV_X80
    CLASS CORE ;
    FOREIGN INV_X80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.840 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.170 0.150 4.95 1.255 ;
        RECT 3.750 0.150 5.375 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.890 0.340 3.06 0.405 ;
        END
    END a
END INV_X80

MACRO INV_Y1
    CLASS CORE ;
    FOREIGN INV_Y1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.760 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.465 0.150 0.53 1.255 ;
        RECT 0.415 0.150 0.61 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.210 0.340 0.34 0.405 ;
        END
    END a
END INV_Y1

MACRO INV_Y2
    CLASS CORE ;
    FOREIGN INV_Y2 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.520 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.925 0.150 1.12 1.255 ;
        RECT 0.835 0.150 1.225 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.420 0.340 0.68 0.405 ;
        END
    END a
END INV_Y2

MACRO INV_Y3
    CLASS CORE ;
    FOREIGN INV_Y3 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.900 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.160 0.150 1.355 1.255 ;
        RECT 1.040 0.150 1.495 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.525 0.340 0.85 0.405 ;
        END
    END a
END INV_Y3

MACRO INV_Y4
    CLASS CORE ;
    FOREIGN INV_Y4 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.900 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.160 0.150 1.355 1.255 ;
        RECT 1.040 0.150 1.495 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.525 0.340 0.85 0.405 ;
        END
    END a
END INV_Y4

MACRO INV_Y6
    CLASS CORE ;
    FOREIGN INV_Y6 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.280 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.150 1.65 1.255 ;
        RECT 1.250 0.150 1.77 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.630 0.340 1.02 0.405 ;
        END
    END a
END INV_Y6

MACRO INV_Y8
    CLASS CORE ;
    FOREIGN INV_Y8 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.620 0.150 1.945 1.255 ;
        RECT 1.460 0.150 2.11 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.735 0.340 1.19 0.405 ;
        END
    END a
END INV_Y8

MACRO INV_Y10
    CLASS CORE ;
    FOREIGN INV_Y10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.620 0.150 1.945 1.255 ;
        RECT 1.460 0.150 2.11 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.735 0.340 1.19 0.405 ;
        END
    END a
END INV_Y10

MACRO INV_Y20
    CLASS CORE ;
    FOREIGN INV_Y20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.315 0.150 2.77 1.255 ;
        RECT 2.085 0.150 2.995 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.050 0.340 1.7 0.405 ;
        END
    END a
END INV_Y20

MACRO INV_Y40
    CLASS CORE ;
    FOREIGN INV_Y40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.940 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.010 0.150 3.595 1.255 ;
        RECT 2.710 0.150 3.88 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.365 0.340 2.21 0.405 ;
        END
    END a
END INV_Y40

MACRO INV_Y80
    CLASS CORE ;
    FOREIGN INV_Y80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.840 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.170 0.150 4.95 1.255 ;
        RECT 3.750 0.150 5.375 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.890 0.340 3.06 0.405 ;
        END
    END a
END INV_Y80

MACRO INV_Z1
    CLASS CORE ;
    FOREIGN INV_Z1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.760 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.465 0.150 0.53 1.255 ;
        RECT 0.415 0.150 0.61 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.210 0.340 0.34 0.405 ;
        END
    END a
END INV_Z1

MACRO INV_Z2
    CLASS CORE ;
    FOREIGN INV_Z2 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.520 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.925 0.150 1.12 1.255 ;
        RECT 0.835 0.150 1.225 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.420 0.340 0.68 0.405 ;
        END
    END a
END INV_Z2

MACRO INV_Z3
    CLASS CORE ;
    FOREIGN INV_Z3 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.900 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.160 0.150 1.355 1.255 ;
        RECT 1.040 0.150 1.495 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.525 0.340 0.85 0.405 ;
        END
    END a
END INV_Z3

MACRO INV_Z4
    CLASS CORE ;
    FOREIGN INV_Z4 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.900 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.160 0.150 1.355 1.255 ;
        RECT 1.040 0.150 1.495 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.525 0.340 0.85 0.405 ;
        END
    END a
END INV_Z4

MACRO INV_Z6
    CLASS CORE ;
    FOREIGN INV_Z6 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.280 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.150 1.65 1.255 ;
        RECT 1.250 0.150 1.77 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.630 0.340 1.02 0.405 ;
        END
    END a
END INV_Z6

MACRO INV_Z8
    CLASS CORE ;
    FOREIGN INV_Z8 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.620 0.150 1.945 1.255 ;
        RECT 1.460 0.150 2.11 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.735 0.340 1.19 0.405 ;
        END
    END a
END INV_Z8

MACRO INV_Z10
    CLASS CORE ;
    FOREIGN INV_Z10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.620 0.150 1.945 1.255 ;
        RECT 1.460 0.150 2.11 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.735 0.340 1.19 0.405 ;
        END
    END a
END INV_Z10

MACRO INV_Z20
    CLASS CORE ;
    FOREIGN INV_Z20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.315 0.150 2.77 1.255 ;
        RECT 2.085 0.150 2.995 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.050 0.340 1.7 0.405 ;
        END
    END a
END INV_Z20

MACRO INV_Z40
    CLASS CORE ;
    FOREIGN INV_Z40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.940 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.010 0.150 3.595 1.255 ;
        RECT 2.710 0.150 3.88 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.365 0.340 2.21 0.405 ;
        END
    END a
END INV_Z40

MACRO INV_Z80
    CLASS CORE ;
    FOREIGN INV_Z80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.840 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.170 0.150 4.95 1.255 ;
        RECT 3.750 0.150 5.375 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.890 0.340 3.06 0.405 ;
        END
    END a
END INV_Z80

MACRO NAND2_X1
    CLASS CORE ;
    FOREIGN NAND2_X1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.140 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.450 0.110 0.58 1.215 ;
        RECT 0.430 0.725 0.625 1.245 ;
        RECT 0.450 0.110 0.905 0.175 ;
        RECT 0.805 0.110 0.935 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.070 0.535 0.33 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.645 0.540 0.905 0.67 ;
        END
    END b
END NAND2_X1

MACRO NAND2_X2
    CLASS CORE ;
    FOREIGN NAND2_X2 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.050 0.110 1.31 1.215 ;
        RECT 1.000 0.725 1.455 1.245 ;
        RECT 1.050 0.110 2.09 0.175 ;
        RECT 1.875 0.110 2.135 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.160 0.535 0.81 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.505 0.540 2.09 0.67 ;
        END
    END b
END NAND2_X2

MACRO NAND2_X3
    CLASS CORE ;
    FOREIGN NAND2_X3 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.420 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.350 0.110 1.675 1.215 ;
        RECT 1.285 0.725 1.87 1.245 ;
        RECT 1.350 0.110 2.715 0.175 ;
        RECT 2.410 0.110 2.735 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.205 0.535 1.05 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.935 0.540 2.715 0.67 ;
        END
    END b
END NAND2_X3

MACRO NAND2_X4
    CLASS CORE ;
    FOREIGN NAND2_X4 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.500 0.110 1.825 1.215 ;
        RECT 1.425 0.725 2.075 1.245 ;
        RECT 1.500 0.110 2.995 0.175 ;
        RECT 2.675 0.110 3.0 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.225 0.535 1.2 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.150 0.540 2.995 0.67 ;
        END
    END b
END NAND2_X4

MACRO NAND2_X6
    CLASS CORE ;
    FOREIGN NAND2_X6 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.800 0.110 2.19 1.215 ;
        RECT 1.710 0.725 2.49 1.245 ;
        RECT 1.800 0.110 3.62 0.175 ;
        RECT 3.210 0.110 3.6 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.270 0.535 1.44 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.580 0.540 3.62 0.67 ;
        END
    END b
END NAND2_X6

MACRO NAND2_X8
    CLASS CORE ;
    FOREIGN NAND2_X8 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.940 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.950 0.110 2.405 1.215 ;
        RECT 1.855 0.725 2.7 1.245 ;
        RECT 1.950 0.110 3.9 0.175 ;
        RECT 3.480 0.110 3.935 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.290 0.535 1.525 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.795 0.540 3.9 0.67 ;
        END
    END b
END NAND2_X8

MACRO NAND2_X10
    CLASS CORE ;
    FOREIGN NAND2_X10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.700 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.250 0.110 2.77 1.215 ;
        RECT 2.140 0.725 3.18 1.245 ;
        RECT 2.250 0.110 4.525 0.175 ;
        RECT 4.015 0.110 4.535 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.340 0.535 1.77 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.225 0.540 4.525 0.67 ;
        END
    END b
END NAND2_X10

MACRO NAND2_X20
    CLASS CORE ;
    FOREIGN NAND2_X20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.000 0.110 3.65 1.215 ;
        RECT 2.850 0.725 4.215 1.245 ;
        RECT 3.000 0.110 5.99 0.175 ;
        RECT 5.350 0.110 6.0 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.450 0.535 2.335 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.300 0.540 6.055 0.67 ;
        END
    END b
END NAND2_X20

MACRO NAND2_X40
    CLASS CORE ;
    FOREIGN NAND2_X40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.200 0.110 5.11 1.215 ;
        RECT 3.990 0.725 5.875 1.245 ;
        RECT 4.200 0.110 8.425 0.175 ;
        RECT 7.490 0.110 8.4 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.630 0.535 3.295 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.020 0.540 8.425 0.67 ;
        END
    END b
END NAND2_X40

MACRO NAND2_X80
    CLASS CORE ;
    FOREIGN NAND2_X80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.440 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.700 0.110 6.935 1.215 ;
        RECT 5.415 0.725 7.95 1.245 ;
        RECT 5.700 0.110 11.42 0.175 ;
        RECT 10.165 0.110 11.4 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.855 0.535 4.495 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.170 0.540 11.42 0.67 ;
        END
    END b
END NAND2_X80

MACRO NAND2_Y01
    CLASS CORE ;
    FOREIGN NAND2_Y01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.140 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.450 0.110 0.58 1.215 ;
        RECT 0.430 0.725 0.625 1.245 ;
        RECT 0.450 0.110 0.905 0.175 ;
        RECT 0.805 0.110 0.935 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.070 0.535 0.33 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.645 0.540 0.905 0.67 ;
        END
    END b
END NAND2_Y01

MACRO NAND2_Y02
    CLASS CORE ;
    FOREIGN NAND2_Y02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.050 0.110 1.31 1.215 ;
        RECT 1.000 0.725 1.455 1.245 ;
        RECT 1.050 0.110 2.09 0.175 ;
        RECT 1.875 0.110 2.135 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.160 0.535 0.81 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.505 0.540 2.09 0.67 ;
        END
    END b
END NAND2_Y02

MACRO NAND2_Y03
    CLASS CORE ;
    FOREIGN NAND2_Y03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.420 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.350 0.110 1.675 1.215 ;
        RECT 1.285 0.725 1.87 1.245 ;
        RECT 1.350 0.110 2.715 0.175 ;
        RECT 2.410 0.110 2.735 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.205 0.535 1.05 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.935 0.540 2.715 0.67 ;
        END
    END b
END NAND2_Y03

MACRO NAND2_Y04
    CLASS CORE ;
    FOREIGN NAND2_Y04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.500 0.110 1.825 1.215 ;
        RECT 1.425 0.725 2.075 1.245 ;
        RECT 1.500 0.110 2.995 0.175 ;
        RECT 2.675 0.110 3.0 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.225 0.535 1.2 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.150 0.540 2.995 0.67 ;
        END
    END b
END NAND2_Y04

MACRO NAND2_Y06
    CLASS CORE ;
    FOREIGN NAND2_Y06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.800 0.110 2.19 1.215 ;
        RECT 1.710 0.725 2.49 1.245 ;
        RECT 1.800 0.110 3.62 0.175 ;
        RECT 3.210 0.110 3.6 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.270 0.535 1.44 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.580 0.540 3.62 0.67 ;
        END
    END b
END NAND2_Y06

MACRO NAND2_Y08
    CLASS CORE ;
    FOREIGN NAND2_Y08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.940 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.950 0.110 2.405 1.215 ;
        RECT 1.855 0.725 2.7 1.245 ;
        RECT 1.950 0.110 3.9 0.175 ;
        RECT 3.480 0.110 3.935 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.290 0.535 1.525 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.795 0.540 3.9 0.67 ;
        END
    END b
END NAND2_Y08

MACRO NAND2_Y10
    CLASS CORE ;
    FOREIGN NAND2_Y10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.700 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.250 0.110 2.77 1.215 ;
        RECT 2.140 0.725 3.18 1.245 ;
        RECT 2.250 0.110 4.525 0.175 ;
        RECT 4.015 0.110 4.535 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.340 0.535 1.77 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.225 0.540 4.525 0.67 ;
        END
    END b
END NAND2_Y10

MACRO NAND2_Y20
    CLASS CORE ;
    FOREIGN NAND2_Y20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.000 0.110 3.65 1.215 ;
        RECT 2.850 0.725 4.215 1.245 ;
        RECT 3.000 0.110 5.99 0.175 ;
        RECT 5.350 0.110 6.0 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.450 0.535 2.335 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.300 0.540 6.055 0.67 ;
        END
    END b
END NAND2_Y20

MACRO NAND2_Y40
    CLASS CORE ;
    FOREIGN NAND2_Y40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.200 0.110 5.11 1.215 ;
        RECT 3.990 0.725 5.875 1.245 ;
        RECT 4.200 0.110 8.425 0.175 ;
        RECT 7.490 0.110 8.4 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.630 0.535 3.295 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.020 0.540 8.425 0.67 ;
        END
    END b
END NAND2_Y40

MACRO NAND2_Y80
    CLASS CORE ;
    FOREIGN NAND2_Y80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.440 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.700 0.110 6.935 1.215 ;
        RECT 5.415 0.725 7.95 1.245 ;
        RECT 5.700 0.110 11.42 0.175 ;
        RECT 10.165 0.110 11.4 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.855 0.535 4.495 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.170 0.540 11.42 0.67 ;
        END
    END b
END NAND2_Y80

MACRO NAND2_Z01
    CLASS CORE ;
    FOREIGN NAND2_Z01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.140 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.450 0.110 0.58 1.215 ;
        RECT 0.430 0.725 0.625 1.245 ;
        RECT 0.450 0.110 0.905 0.175 ;
        RECT 0.805 0.110 0.935 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.070 0.535 0.33 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.645 0.540 0.905 0.67 ;
        END
    END b
END NAND2_Z01

MACRO NAND2_Z02
    CLASS CORE ;
    FOREIGN NAND2_Z02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.050 0.110 1.31 1.215 ;
        RECT 1.000 0.725 1.455 1.245 ;
        RECT 1.050 0.110 2.09 0.175 ;
        RECT 1.875 0.110 2.135 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.160 0.535 0.81 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.505 0.540 2.09 0.67 ;
        END
    END b
END NAND2_Z02

MACRO NAND2_Z03
    CLASS CORE ;
    FOREIGN NAND2_Z03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.420 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.350 0.110 1.675 1.215 ;
        RECT 1.285 0.725 1.87 1.245 ;
        RECT 1.350 0.110 2.715 0.175 ;
        RECT 2.410 0.110 2.735 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.205 0.535 1.05 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.935 0.540 2.715 0.67 ;
        END
    END b
END NAND2_Z03

MACRO NAND2_Z04
    CLASS CORE ;
    FOREIGN NAND2_Z04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.500 0.110 1.825 1.215 ;
        RECT 1.425 0.725 2.075 1.245 ;
        RECT 1.500 0.110 2.995 0.175 ;
        RECT 2.675 0.110 3.0 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.225 0.535 1.2 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.150 0.540 2.995 0.67 ;
        END
    END b
END NAND2_Z04

MACRO NAND2_Z06
    CLASS CORE ;
    FOREIGN NAND2_Z06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.800 0.110 2.19 1.215 ;
        RECT 1.710 0.725 2.49 1.245 ;
        RECT 1.800 0.110 3.62 0.175 ;
        RECT 3.210 0.110 3.6 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.270 0.535 1.44 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.580 0.540 3.62 0.67 ;
        END
    END b
END NAND2_Z06

MACRO NAND2_Z08
    CLASS CORE ;
    FOREIGN NAND2_Z08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.940 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.950 0.110 2.405 1.215 ;
        RECT 1.855 0.725 2.7 1.245 ;
        RECT 1.950 0.110 3.9 0.175 ;
        RECT 3.480 0.110 3.935 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.290 0.535 1.525 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.795 0.540 3.9 0.67 ;
        END
    END b
END NAND2_Z08

MACRO NAND2_Z10
    CLASS CORE ;
    FOREIGN NAND2_Z10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.700 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.250 0.110 2.77 1.215 ;
        RECT 2.140 0.725 3.18 1.245 ;
        RECT 2.250 0.110 4.525 0.175 ;
        RECT 4.015 0.110 4.535 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.340 0.535 1.77 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.225 0.540 4.525 0.67 ;
        END
    END b
END NAND2_Z10

MACRO NAND2_Z20
    CLASS CORE ;
    FOREIGN NAND2_Z20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.000 0.110 3.65 1.215 ;
        RECT 2.850 0.725 4.215 1.245 ;
        RECT 3.000 0.110 5.99 0.175 ;
        RECT 5.350 0.110 6.0 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.450 0.535 2.335 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.300 0.540 6.055 0.67 ;
        END
    END b
END NAND2_Z20

MACRO NAND2_Z40
    CLASS CORE ;
    FOREIGN NAND2_Z40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.200 0.110 5.11 1.215 ;
        RECT 3.990 0.725 5.875 1.245 ;
        RECT 4.200 0.110 8.425 0.175 ;
        RECT 7.490 0.110 8.4 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.630 0.535 3.295 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.020 0.540 8.425 0.67 ;
        END
    END b
END NAND2_Z40

MACRO NAND2_Z80
    CLASS CORE ;
    FOREIGN NAND2_Z80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.440 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.700 0.110 6.935 1.215 ;
        RECT 5.415 0.725 7.95 1.245 ;
        RECT 5.700 0.110 11.42 0.175 ;
        RECT 10.165 0.110 11.4 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.855 0.535 4.495 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.170 0.540 11.42 0.67 ;
        END
    END b
END NAND2_Z80

MACRO NAND3_X1
    CLASS CORE ;
    FOREIGN NAND3_X1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.140 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.415 0.805 0.48 1.26 ;
        RECT 0.415 0.805 0.935 0.87 ;
        RECT 0.875 0.090 0.94 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.040 0.630 0.3 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.350 0.090 0.545 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.640 0.090 0.77 0.74 ;
        END
    END c
END NAND3_X1

MACRO NAND3_X2
    CLASS CORE ;
    FOREIGN NAND3_X2 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.975 0.805 1.17 1.26 ;
        RECT 0.975 0.805 2.21 0.87 ;
        RECT 2.035 0.090 2.23 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.090 0.630 0.61 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.820 0.090 1.34 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.490 0.090 1.815 0.74 ;
        END
    END c
END NAND3_X2

MACRO NAND3_X3
    CLASS CORE ;
    FOREIGN NAND3_X3 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.420 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.250 0.805 1.51 1.26 ;
        RECT 1.250 0.805 2.875 0.87 ;
        RECT 2.620 0.090 2.88 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.115 0.630 0.83 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.055 0.090 1.705 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.915 0.090 2.37 0.74 ;
        END
    END c
END NAND3_X3

MACRO NAND3_X4
    CLASS CORE ;
    FOREIGN NAND3_X4 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.805 1.65 1.26 ;
        RECT 1.390 0.805 3.145 0.87 ;
        RECT 2.910 0.090 3.17 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.130 0.630 0.91 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.170 0.090 1.885 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.130 0.090 2.65 0.74 ;
        END
    END c
END NAND3_X4

MACRO NAND3_X6
    CLASS CORE ;
    FOREIGN NAND3_X6 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.670 0.805 1.995 1.26 ;
        RECT 1.670 0.805 3.815 0.87 ;
        RECT 3.490 0.090 3.815 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.155 0.630 1.065 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.405 0.090 2.25 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.555 0.090 3.14 0.74 ;
        END
    END c
END NAND3_X6

MACRO NAND3_X8
    CLASS CORE ;
    FOREIGN NAND3_X8 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.940 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.805 0.805 2.13 1.26 ;
        RECT 1.805 0.805 4.145 0.87 ;
        RECT 3.785 0.090 4.11 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.170 0.630 1.145 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.520 0.090 2.43 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.770 0.090 3.42 0.74 ;
        END
    END c
END NAND3_X8

MACRO NAND3_X10
    CLASS CORE ;
    FOREIGN NAND3_X10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.700 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.085 0.805 2.475 1.26 ;
        RECT 2.085 0.805 4.75 0.87 ;
        RECT 4.365 0.090 4.755 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.195 0.630 1.365 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.755 0.090 2.795 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.195 0.090 3.975 0.74 ;
        END
    END c
END NAND3_X10

MACRO NAND3_X20
    CLASS CORE ;
    FOREIGN NAND3_X20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.780 0.805 3.3 1.26 ;
        RECT 2.780 0.805 6.355 0.87 ;
        RECT 5.820 0.090 6.34 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.260 0.630 1.755 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.340 0.090 3.77 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.260 0.090 5.235 0.74 ;
        END
    END c
END NAND3_X20

MACRO NAND3_X40
    CLASS CORE ;
    FOREIGN NAND3_X40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.890 0.805 4.605 1.26 ;
        RECT 3.890 0.805 8.895 0.87 ;
        RECT 8.150 0.090 8.865 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.365 0.630 2.51 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.275 0.090 5.225 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.965 0.090 7.395 0.74 ;
        END
    END c
END NAND3_X40

MACRO NAND3_X80
    CLASS CORE ;
    FOREIGN NAND3_X80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.440 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.280 0.805 6.255 1.26 ;
        RECT 5.280 0.805 12.04 0.87 ;
        RECT 11.060 0.090 12.035 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.495 0.630 3.355 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.445 0.090 7.11 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.095 0.090 9.98 0.74 ;
        END
    END c
END NAND3_X80

MACRO NAND3_Y1
    CLASS CORE ;
    FOREIGN NAND3_Y1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.140 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.415 0.805 0.48 1.26 ;
        RECT 0.415 0.805 0.935 0.87 ;
        RECT 0.875 0.090 0.94 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.040 0.630 0.3 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.350 0.090 0.545 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.640 0.090 0.77 0.74 ;
        END
    END c
END NAND3_Y1

MACRO NAND3_Y2
    CLASS CORE ;
    FOREIGN NAND3_Y2 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.975 0.805 1.17 1.26 ;
        RECT 0.975 0.805 2.21 0.87 ;
        RECT 2.035 0.090 2.23 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.090 0.630 0.61 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.820 0.090 1.34 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.490 0.090 1.815 0.74 ;
        END
    END c
END NAND3_Y2

MACRO NAND3_Y3
    CLASS CORE ;
    FOREIGN NAND3_Y3 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.420 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.250 0.805 1.51 1.26 ;
        RECT 1.250 0.805 2.875 0.87 ;
        RECT 2.620 0.090 2.88 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.115 0.630 0.83 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.055 0.090 1.705 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.915 0.090 2.37 0.74 ;
        END
    END c
END NAND3_Y3

MACRO NAND3_Y4
    CLASS CORE ;
    FOREIGN NAND3_Y4 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.805 1.65 1.26 ;
        RECT 1.390 0.805 3.145 0.87 ;
        RECT 2.910 0.090 3.17 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.130 0.630 0.91 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.170 0.090 1.885 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.130 0.090 2.65 0.74 ;
        END
    END c
END NAND3_Y4

MACRO NAND3_Y6
    CLASS CORE ;
    FOREIGN NAND3_Y6 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.670 0.805 1.995 1.26 ;
        RECT 1.670 0.805 3.815 0.87 ;
        RECT 3.490 0.090 3.815 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.155 0.630 1.065 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.405 0.090 2.25 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.555 0.090 3.14 0.74 ;
        END
    END c
END NAND3_Y6

MACRO NAND3_Y8
    CLASS CORE ;
    FOREIGN NAND3_Y8 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.940 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.805 0.805 2.13 1.26 ;
        RECT 1.805 0.805 4.145 0.87 ;
        RECT 3.785 0.090 4.11 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.170 0.630 1.145 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.520 0.090 2.43 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.770 0.090 3.42 0.74 ;
        END
    END c
END NAND3_Y8

MACRO NAND3_Y10
    CLASS CORE ;
    FOREIGN NAND3_Y10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.700 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.085 0.805 2.475 1.26 ;
        RECT 2.085 0.805 4.75 0.87 ;
        RECT 4.365 0.090 4.755 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.195 0.630 1.365 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.755 0.090 2.795 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.195 0.090 3.975 0.74 ;
        END
    END c
END NAND3_Y10

MACRO NAND3_Y20
    CLASS CORE ;
    FOREIGN NAND3_Y20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.780 0.805 3.3 1.26 ;
        RECT 2.780 0.805 6.355 0.87 ;
        RECT 5.820 0.090 6.34 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.260 0.630 1.755 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.340 0.090 3.77 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.260 0.090 5.235 0.74 ;
        END
    END c
END NAND3_Y20

MACRO NAND3_Y40
    CLASS CORE ;
    FOREIGN NAND3_Y40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.890 0.805 4.605 1.26 ;
        RECT 3.890 0.805 8.895 0.87 ;
        RECT 8.150 0.090 8.865 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.365 0.630 2.51 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.275 0.090 5.225 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.965 0.090 7.395 0.74 ;
        END
    END c
END NAND3_Y40

MACRO NAND3_Y80
    CLASS CORE ;
    FOREIGN NAND3_Y80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.440 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.280 0.805 6.255 1.26 ;
        RECT 5.280 0.805 12.04 0.87 ;
        RECT 11.060 0.090 12.035 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.495 0.630 3.355 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.445 0.090 7.11 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.095 0.090 9.98 0.74 ;
        END
    END c
END NAND3_Y80

MACRO NAND3_Z1
    CLASS CORE ;
    FOREIGN NAND3_Z1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.140 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.415 0.805 0.48 1.26 ;
        RECT 0.415 0.805 0.935 0.87 ;
        RECT 0.875 0.090 0.94 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.040 0.630 0.3 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.350 0.090 0.545 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.640 0.090 0.77 0.74 ;
        END
    END c
END NAND3_Z1

MACRO NAND3_Z2
    CLASS CORE ;
    FOREIGN NAND3_Z2 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.975 0.805 1.17 1.26 ;
        RECT 0.975 0.805 2.21 0.87 ;
        RECT 2.035 0.090 2.23 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.090 0.630 0.61 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.820 0.090 1.34 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.490 0.090 1.815 0.74 ;
        END
    END c
END NAND3_Z2

MACRO NAND3_Z3
    CLASS CORE ;
    FOREIGN NAND3_Z3 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.420 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.250 0.805 1.51 1.26 ;
        RECT 1.250 0.805 2.875 0.87 ;
        RECT 2.620 0.090 2.88 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.115 0.630 0.83 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.055 0.090 1.705 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.915 0.090 2.37 0.74 ;
        END
    END c
END NAND3_Z3

MACRO NAND3_Z4
    CLASS CORE ;
    FOREIGN NAND3_Z4 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.805 1.65 1.26 ;
        RECT 1.390 0.805 3.145 0.87 ;
        RECT 2.910 0.090 3.17 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.130 0.630 0.91 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.170 0.090 1.885 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.130 0.090 2.65 0.74 ;
        END
    END c
END NAND3_Z4

MACRO NAND3_Z6
    CLASS CORE ;
    FOREIGN NAND3_Z6 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.670 0.805 1.995 1.26 ;
        RECT 1.670 0.805 3.815 0.87 ;
        RECT 3.490 0.090 3.815 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.155 0.630 1.065 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.405 0.090 2.25 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.555 0.090 3.14 0.74 ;
        END
    END c
END NAND3_Z6

MACRO NAND3_Z8
    CLASS CORE ;
    FOREIGN NAND3_Z8 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.940 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.805 0.805 2.13 1.26 ;
        RECT 1.805 0.805 4.145 0.87 ;
        RECT 3.785 0.090 4.11 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.170 0.630 1.145 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.520 0.090 2.43 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.770 0.090 3.42 0.74 ;
        END
    END c
END NAND3_Z8

MACRO NAND3_Z10
    CLASS CORE ;
    FOREIGN NAND3_Z10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.700 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.085 0.805 2.475 1.26 ;
        RECT 2.085 0.805 4.75 0.87 ;
        RECT 4.365 0.090 4.755 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.195 0.630 1.365 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.755 0.090 2.795 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.195 0.090 3.975 0.74 ;
        END
    END c
END NAND3_Z10

MACRO NAND3_Z20
    CLASS CORE ;
    FOREIGN NAND3_Z20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.780 0.805 3.3 1.26 ;
        RECT 2.780 0.805 6.355 0.87 ;
        RECT 5.820 0.090 6.34 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.260 0.630 1.755 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.340 0.090 3.77 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.260 0.090 5.235 0.74 ;
        END
    END c
END NAND3_Z20

MACRO NAND3_Z40
    CLASS CORE ;
    FOREIGN NAND3_Z40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.890 0.805 4.605 1.26 ;
        RECT 3.890 0.805 8.895 0.87 ;
        RECT 8.150 0.090 8.865 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.365 0.630 2.51 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.275 0.090 5.225 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.965 0.090 7.395 0.74 ;
        END
    END c
END NAND3_Z40

MACRO NAND3_Z80
    CLASS CORE ;
    FOREIGN NAND3_Z80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.440 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.280 0.805 6.255 1.26 ;
        RECT 5.280 0.805 12.04 0.87 ;
        RECT 11.060 0.090 12.035 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.495 0.630 3.355 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.445 0.090 7.11 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.095 0.090 9.98 0.74 ;
        END
    END c
END NAND3_Z80

MACRO NAND4_X1
    CLASS CORE ;
    FOREIGN NAND4_X1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.520 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.465 0.210 0.53 0.925 ;
        RECT 0.465 0.870 0.79 0.935 ;
        RECT 0.715 0.870 0.78 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.145 0.725 1.34 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.890 0.725 1.085 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.210 0.635 0.405 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.635 0.725 0.83 0.79 ;
        END
    END d
END NAND4_X1

MACRO NAND4_X2
    CLASS CORE ;
    FOREIGN NAND4_X2 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.040 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.925 0.210 1.12 0.925 ;
        RECT 0.925 0.870 1.575 0.935 ;
        RECT 1.435 0.870 1.63 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.285 0.725 2.61 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.780 0.725 2.105 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.420 0.635 0.745 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.275 0.725 1.6 0.79 ;
        END
    END d
END NAND4_X2

MACRO NAND4_X3
    CLASS CORE ;
    FOREIGN NAND4_X3 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.160 0.210 1.355 0.925 ;
        RECT 1.160 0.870 2.005 0.935 ;
        RECT 1.790 0.870 1.985 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.860 0.725 3.25 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.225 0.725 2.615 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.525 0.635 0.915 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.590 0.725 1.98 0.79 ;
        END
    END d
END NAND4_X3

MACRO NAND4_X4
    CLASS CORE ;
    FOREIGN NAND4_X4 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.210 1.65 0.925 ;
        RECT 1.390 0.870 2.43 0.935 ;
        RECT 2.150 0.870 2.41 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.430 0.725 3.95 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.670 0.725 3.19 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.630 0.635 1.15 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.910 0.725 2.43 0.79 ;
        END
    END d
END NAND4_X4

MACRO NAND4_X6
    CLASS CORE ;
    FOREIGN NAND4_X6 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.620 0.210 1.945 0.925 ;
        RECT 1.620 0.870 2.79 0.935 ;
        RECT 2.510 0.870 2.835 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.000 0.725 4.585 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.115 0.725 3.7 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.735 0.635 1.32 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.230 0.725 2.815 0.79 ;
        END
    END d
END NAND4_X6

MACRO NAND4_X8
    CLASS CORE ;
    FOREIGN NAND4_X8 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.080 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.855 0.210 2.18 0.925 ;
        RECT 1.855 0.870 3.22 0.935 ;
        RECT 2.865 0.870 3.19 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.575 0.725 5.225 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.560 0.725 4.21 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.840 0.635 1.49 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.545 0.725 3.195 0.79 ;
        END
    END d
END NAND4_X8

MACRO NAND4_X10
    CLASS CORE ;
    FOREIGN NAND4_X10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.460 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.970 0.210 2.36 0.925 ;
        RECT 1.970 0.870 3.4 0.935 ;
        RECT 3.045 0.870 3.435 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.860 0.725 5.575 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.785 0.725 4.5 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.895 0.635 1.61 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.705 0.725 3.42 0.79 ;
        END
    END d
END NAND4_X10

MACRO NAND4_X20
    CLASS CORE ;
    FOREIGN NAND4_X20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.740 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.665 0.210 3.185 0.925 ;
        RECT 2.665 0.870 4.615 0.935 ;
        RECT 4.120 0.870 4.64 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.575 0.725 7.55 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.115 0.725 6.09 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.210 0.635 2.185 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.660 0.725 4.635 0.79 ;
        END
    END d
END NAND4_X20

MACRO NAND4_X40
    CLASS CORE ;
    FOREIGN NAND4_X40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.780 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.590 0.210 4.24 0.925 ;
        RECT 3.590 0.870 6.255 0.935 ;
        RECT 5.555 0.870 6.205 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.860 0.725 10.16 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.895 0.725 8.195 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.625 0.635 2.925 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.935 0.725 6.235 0.79 ;
        END
    END d
END NAND4_X40

MACRO NAND4_X80
    CLASS CORE ;
    FOREIGN NAND4_X80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.340 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.980 0.210 5.89 0.925 ;
        RECT 4.980 0.870 8.62 0.935 ;
        RECT 7.705 0.870 8.615 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 12.290 0.725 14.11 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 9.565 0.725 11.385 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.255 0.635 4.075 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.845 0.725 8.665 0.79 ;
        END
    END d
END NAND4_X80

MACRO NAND4_Y1
    CLASS CORE ;
    FOREIGN NAND4_Y1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.520 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.465 0.210 0.53 0.925 ;
        RECT 0.465 0.870 0.79 0.935 ;
        RECT 0.715 0.870 0.78 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.145 0.725 1.34 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.890 0.725 1.085 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.210 0.635 0.405 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.635 0.725 0.83 0.79 ;
        END
    END d
END NAND4_Y1

MACRO NAND4_Y2
    CLASS CORE ;
    FOREIGN NAND4_Y2 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.040 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.925 0.210 1.12 0.925 ;
        RECT 0.925 0.870 1.575 0.935 ;
        RECT 1.435 0.870 1.63 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.285 0.725 2.61 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.780 0.725 2.105 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.420 0.635 0.745 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.275 0.725 1.6 0.79 ;
        END
    END d
END NAND4_Y2

MACRO NAND4_Y3
    CLASS CORE ;
    FOREIGN NAND4_Y3 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.160 0.210 1.355 0.925 ;
        RECT 1.160 0.870 2.005 0.935 ;
        RECT 1.790 0.870 1.985 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.860 0.725 3.25 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.225 0.725 2.615 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.525 0.635 0.915 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.590 0.725 1.98 0.79 ;
        END
    END d
END NAND4_Y3

MACRO NAND4_Y4
    CLASS CORE ;
    FOREIGN NAND4_Y4 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.210 1.65 0.925 ;
        RECT 1.390 0.870 2.43 0.935 ;
        RECT 2.150 0.870 2.41 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.430 0.725 3.95 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.670 0.725 3.19 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.630 0.635 1.15 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.910 0.725 2.43 0.79 ;
        END
    END d
END NAND4_Y4

MACRO NAND4_Y6
    CLASS CORE ;
    FOREIGN NAND4_Y6 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.620 0.210 1.945 0.925 ;
        RECT 1.620 0.870 2.79 0.935 ;
        RECT 2.510 0.870 2.835 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.000 0.725 4.585 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.115 0.725 3.7 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.735 0.635 1.32 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.230 0.725 2.815 0.79 ;
        END
    END d
END NAND4_Y6

MACRO NAND4_Y8
    CLASS CORE ;
    FOREIGN NAND4_Y8 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.080 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.855 0.210 2.18 0.925 ;
        RECT 1.855 0.870 3.22 0.935 ;
        RECT 2.865 0.870 3.19 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.575 0.725 5.225 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.560 0.725 4.21 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.840 0.635 1.49 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.545 0.725 3.195 0.79 ;
        END
    END d
END NAND4_Y8

MACRO NAND4_Y10
    CLASS CORE ;
    FOREIGN NAND4_Y10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.460 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.970 0.210 2.36 0.925 ;
        RECT 1.970 0.870 3.4 0.935 ;
        RECT 3.045 0.870 3.435 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.860 0.725 5.575 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.785 0.725 4.5 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.895 0.635 1.61 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.705 0.725 3.42 0.79 ;
        END
    END d
END NAND4_Y10

MACRO NAND4_Y20
    CLASS CORE ;
    FOREIGN NAND4_Y20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.740 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.665 0.210 3.185 0.925 ;
        RECT 2.665 0.870 4.615 0.935 ;
        RECT 4.120 0.870 4.64 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.575 0.725 7.55 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.115 0.725 6.09 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.210 0.635 2.185 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.660 0.725 4.635 0.79 ;
        END
    END d
END NAND4_Y20

MACRO NAND4_Y40
    CLASS CORE ;
    FOREIGN NAND4_Y40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.780 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.590 0.210 4.24 0.925 ;
        RECT 3.590 0.870 6.255 0.935 ;
        RECT 5.555 0.870 6.205 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.860 0.725 10.16 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.895 0.725 8.195 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.625 0.635 2.925 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.935 0.725 6.235 0.79 ;
        END
    END d
END NAND4_Y40

MACRO NAND4_Y80
    CLASS CORE ;
    FOREIGN NAND4_Y80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.340 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.980 0.210 5.89 0.925 ;
        RECT 4.980 0.870 8.62 0.935 ;
        RECT 7.705 0.870 8.615 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 12.290 0.725 14.11 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 9.565 0.725 11.385 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.255 0.635 4.075 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.845 0.725 8.665 0.79 ;
        END
    END d
END NAND4_Y80

MACRO NAND4_Z1
    CLASS CORE ;
    FOREIGN NAND4_Z1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.520 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.465 0.210 0.53 0.925 ;
        RECT 0.465 0.870 0.79 0.935 ;
        RECT 0.715 0.870 0.78 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.145 0.725 1.34 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.890 0.725 1.085 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.210 0.635 0.405 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.635 0.725 0.83 0.79 ;
        END
    END d
END NAND4_Z1

MACRO NAND4_Z2
    CLASS CORE ;
    FOREIGN NAND4_Z2 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.040 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.925 0.210 1.12 0.925 ;
        RECT 0.925 0.870 1.575 0.935 ;
        RECT 1.435 0.870 1.63 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.285 0.725 2.61 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.780 0.725 2.105 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.420 0.635 0.745 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.275 0.725 1.6 0.79 ;
        END
    END d
END NAND4_Z2

MACRO NAND4_Z3
    CLASS CORE ;
    FOREIGN NAND4_Z3 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.160 0.210 1.355 0.925 ;
        RECT 1.160 0.870 2.005 0.935 ;
        RECT 1.790 0.870 1.985 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.860 0.725 3.25 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.225 0.725 2.615 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.525 0.635 0.915 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.590 0.725 1.98 0.79 ;
        END
    END d
END NAND4_Z3

MACRO NAND4_Z4
    CLASS CORE ;
    FOREIGN NAND4_Z4 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.210 1.65 0.925 ;
        RECT 1.390 0.870 2.43 0.935 ;
        RECT 2.150 0.870 2.41 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.430 0.725 3.95 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.670 0.725 3.19 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.630 0.635 1.15 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.910 0.725 2.43 0.79 ;
        END
    END d
END NAND4_Z4

MACRO NAND4_Z6
    CLASS CORE ;
    FOREIGN NAND4_Z6 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.620 0.210 1.945 0.925 ;
        RECT 1.620 0.870 2.79 0.935 ;
        RECT 2.510 0.870 2.835 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.000 0.725 4.585 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.115 0.725 3.7 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.735 0.635 1.32 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.230 0.725 2.815 0.79 ;
        END
    END d
END NAND4_Z6

MACRO NAND4_Z8
    CLASS CORE ;
    FOREIGN NAND4_Z8 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.080 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.855 0.210 2.18 0.925 ;
        RECT 1.855 0.870 3.22 0.935 ;
        RECT 2.865 0.870 3.19 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.575 0.725 5.225 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.560 0.725 4.21 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.840 0.635 1.49 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.545 0.725 3.195 0.79 ;
        END
    END d
END NAND4_Z8

MACRO NAND4_Z10
    CLASS CORE ;
    FOREIGN NAND4_Z10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.460 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.970 0.210 2.36 0.925 ;
        RECT 1.970 0.870 3.4 0.935 ;
        RECT 3.045 0.870 3.435 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.860 0.725 5.575 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.785 0.725 4.5 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.895 0.635 1.61 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.705 0.725 3.42 0.79 ;
        END
    END d
END NAND4_Z10

MACRO NAND4_Z20
    CLASS CORE ;
    FOREIGN NAND4_Z20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.740 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.665 0.210 3.185 0.925 ;
        RECT 2.665 0.870 4.615 0.935 ;
        RECT 4.120 0.870 4.64 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.575 0.725 7.55 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.115 0.725 6.09 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.210 0.635 2.185 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.660 0.725 4.635 0.79 ;
        END
    END d
END NAND4_Z20

MACRO NAND4_Z40
    CLASS CORE ;
    FOREIGN NAND4_Z40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.780 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.590 0.210 4.24 0.925 ;
        RECT 3.590 0.870 6.255 0.935 ;
        RECT 5.555 0.870 6.205 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.860 0.725 10.16 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.895 0.725 8.195 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.625 0.635 2.925 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.935 0.725 6.235 0.79 ;
        END
    END d
END NAND4_Z40

MACRO NAND4_Z80
    CLASS CORE ;
    FOREIGN NAND4_Z80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.340 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.980 0.210 5.89 0.925 ;
        RECT 4.980 0.870 8.62 0.935 ;
        RECT 7.705 0.870 8.615 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 12.290 0.725 14.11 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 9.565 0.725 11.385 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.255 0.635 4.075 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.845 0.725 8.665 0.79 ;
        END
    END d
END NAND4_Z80

MACRO NOR2_X1
    CLASS CORE ;
    FOREIGN NOR2_X1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.140 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.520 0.150 0.65 0.54 ;
        RECT 0.465 0.150 0.66 0.28 ;
        RECT 0.520 0.505 0.91 0.57 ;
        RECT 0.805 0.505 0.935 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.235 0.340 0.43 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.715 0.340 0.91 0.405 ;
        END
    END b
END NOR2_X1

MACRO NOR2_X2
    CLASS CORE ;
    FOREIGN NOR2_X2 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.215 0.150 1.475 0.54 ;
        RECT 1.085 0.150 1.54 0.28 ;
        RECT 1.215 0.505 2.125 0.57 ;
        RECT 1.875 0.505 2.135 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.550 0.340 1.005 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.670 0.340 2.125 0.405 ;
        END
    END b
END NOR2_X2

MACRO NOR2_X3
    CLASS CORE ;
    FOREIGN NOR2_X3 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.420 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.565 0.150 1.89 0.54 ;
        RECT 1.395 0.150 1.98 0.28 ;
        RECT 1.565 0.505 2.67 0.57 ;
        RECT 2.410 0.505 2.735 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.710 0.340 1.295 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.150 0.340 2.735 0.405 ;
        END
    END b
END NOR2_X3

MACRO NOR2_X4
    CLASS CORE ;
    FOREIGN NOR2_X4 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.740 0.150 2.065 0.54 ;
        RECT 1.550 0.150 2.2 0.28 ;
        RECT 1.740 0.505 2.975 0.57 ;
        RECT 2.675 0.505 3.0 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.790 0.340 1.44 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.390 0.340 3.04 0.405 ;
        END
    END b
END NOR2_X4

MACRO NOR2_X6
    CLASS CORE ;
    FOREIGN NOR2_X6 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.085 0.150 2.475 0.54 ;
        RECT 1.860 0.150 2.64 0.28 ;
        RECT 2.085 0.505 3.58 0.57 ;
        RECT 3.210 0.505 3.6 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.945 0.340 1.725 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.865 0.340 3.645 0.405 ;
        END
    END b
END NOR2_X6

MACRO NOR2_X8
    CLASS CORE ;
    FOREIGN NOR2_X8 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.940 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.260 0.150 2.715 0.54 ;
        RECT 2.015 0.150 2.86 0.28 ;
        RECT 2.260 0.505 3.885 0.57 ;
        RECT 3.480 0.505 3.935 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.025 0.340 1.87 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.105 0.340 3.95 0.405 ;
        END
    END b
END NOR2_X8

MACRO NOR2_X10
    CLASS CORE ;
    FOREIGN NOR2_X10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.700 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.605 0.150 3.125 0.54 ;
        RECT 2.325 0.150 3.365 0.28 ;
        RECT 2.605 0.505 4.49 0.57 ;
        RECT 4.015 0.505 4.535 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.180 0.340 2.09 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.580 0.340 4.49 0.405 ;
        END
    END b
END NOR2_X10

MACRO NOR2_X20
    CLASS CORE ;
    FOREIGN NOR2_X20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.475 0.150 4.125 0.54 ;
        RECT 3.100 0.150 4.465 0.28 ;
        RECT 3.475 0.505 6.01 0.57 ;
        RECT 5.350 0.505 6.0 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.575 0.340 2.81 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.775 0.340 6.01 0.405 ;
        END
    END b
END NOR2_X20

MACRO NOR2_X40
    CLASS CORE ;
    FOREIGN NOR2_X40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.865 0.150 5.775 0.54 ;
        RECT 4.340 0.150 6.225 0.28 ;
        RECT 4.865 0.505 8.375 0.57 ;
        RECT 7.490 0.505 8.4 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.205 0.340 3.96 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.685 0.340 8.44 0.405 ;
        END
    END b
END NOR2_X40

MACRO NOR2_X80
    CLASS CORE ;
    FOREIGN NOR2_X80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.440 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.605 0.150 7.84 0.54 ;
        RECT 5.890 0.150 8.425 0.28 ;
        RECT 6.605 0.505 11.415 0.57 ;
        RECT 10.165 0.505 11.4 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.995 0.340 5.4 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 9.075 0.340 11.48 0.405 ;
        END
    END b
END NOR2_X80

MACRO NOR2_Y1
    CLASS CORE ;
    FOREIGN NOR2_Y1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.140 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.520 0.150 0.65 0.54 ;
        RECT 0.465 0.150 0.66 0.28 ;
        RECT 0.520 0.505 0.91 0.57 ;
        RECT 0.805 0.505 0.935 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.235 0.340 0.43 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.715 0.340 0.91 0.405 ;
        END
    END b
END NOR2_Y1

MACRO NOR2_Y2
    CLASS CORE ;
    FOREIGN NOR2_Y2 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.215 0.150 1.475 0.54 ;
        RECT 1.085 0.150 1.54 0.28 ;
        RECT 1.215 0.505 2.125 0.57 ;
        RECT 1.875 0.505 2.135 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.550 0.340 1.005 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.670 0.340 2.125 0.405 ;
        END
    END b
END NOR2_Y2

MACRO NOR2_Y3
    CLASS CORE ;
    FOREIGN NOR2_Y3 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.420 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.565 0.150 1.89 0.54 ;
        RECT 1.395 0.150 1.98 0.28 ;
        RECT 1.565 0.505 2.67 0.57 ;
        RECT 2.410 0.505 2.735 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.710 0.340 1.295 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.150 0.340 2.735 0.405 ;
        END
    END b
END NOR2_Y3

MACRO NOR2_Y4
    CLASS CORE ;
    FOREIGN NOR2_Y4 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.740 0.150 2.065 0.54 ;
        RECT 1.550 0.150 2.2 0.28 ;
        RECT 1.740 0.505 2.975 0.57 ;
        RECT 2.675 0.505 3.0 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.790 0.340 1.44 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.390 0.340 3.04 0.405 ;
        END
    END b
END NOR2_Y4

MACRO NOR2_Y6
    CLASS CORE ;
    FOREIGN NOR2_Y6 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.085 0.150 2.475 0.54 ;
        RECT 1.860 0.150 2.64 0.28 ;
        RECT 2.085 0.505 3.58 0.57 ;
        RECT 3.210 0.505 3.6 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.945 0.340 1.725 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.865 0.340 3.645 0.405 ;
        END
    END b
END NOR2_Y6

MACRO NOR2_Y8
    CLASS CORE ;
    FOREIGN NOR2_Y8 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.940 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.260 0.150 2.715 0.54 ;
        RECT 2.015 0.150 2.86 0.28 ;
        RECT 2.260 0.505 3.885 0.57 ;
        RECT 3.480 0.505 3.935 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.025 0.340 1.87 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.105 0.340 3.95 0.405 ;
        END
    END b
END NOR2_Y8

MACRO NOR2_Y10
    CLASS CORE ;
    FOREIGN NOR2_Y10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.700 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.605 0.150 3.125 0.54 ;
        RECT 2.325 0.150 3.365 0.28 ;
        RECT 2.605 0.505 4.49 0.57 ;
        RECT 4.015 0.505 4.535 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.180 0.340 2.09 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.580 0.340 4.49 0.405 ;
        END
    END b
END NOR2_Y10

MACRO NOR2_Y20
    CLASS CORE ;
    FOREIGN NOR2_Y20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.475 0.150 4.125 0.54 ;
        RECT 3.100 0.150 4.465 0.28 ;
        RECT 3.475 0.505 6.01 0.57 ;
        RECT 5.350 0.505 6.0 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.575 0.340 2.81 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.775 0.340 6.01 0.405 ;
        END
    END b
END NOR2_Y20

MACRO NOR2_Y40
    CLASS CORE ;
    FOREIGN NOR2_Y40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.865 0.150 5.775 0.54 ;
        RECT 4.340 0.150 6.225 0.28 ;
        RECT 4.865 0.505 8.375 0.57 ;
        RECT 7.490 0.505 8.4 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.205 0.340 3.96 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.685 0.340 8.44 0.405 ;
        END
    END b
END NOR2_Y40

MACRO NOR2_Y80
    CLASS CORE ;
    FOREIGN NOR2_Y80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.440 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.605 0.150 7.84 0.54 ;
        RECT 5.890 0.150 8.425 0.28 ;
        RECT 6.605 0.505 11.415 0.57 ;
        RECT 10.165 0.505 11.4 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.995 0.340 5.4 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 9.075 0.340 11.48 0.405 ;
        END
    END b
END NOR2_Y80

MACRO NOR2_Z1
    CLASS CORE ;
    FOREIGN NOR2_Z1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.140 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.520 0.150 0.65 0.54 ;
        RECT 0.465 0.150 0.66 0.28 ;
        RECT 0.520 0.505 0.91 0.57 ;
        RECT 0.805 0.505 0.935 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.235 0.340 0.43 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.715 0.340 0.91 0.405 ;
        END
    END b
END NOR2_Z1

MACRO NOR2_Z2
    CLASS CORE ;
    FOREIGN NOR2_Z2 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.215 0.150 1.475 0.54 ;
        RECT 1.085 0.150 1.54 0.28 ;
        RECT 1.215 0.505 2.125 0.57 ;
        RECT 1.875 0.505 2.135 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.550 0.340 1.005 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.670 0.340 2.125 0.405 ;
        END
    END b
END NOR2_Z2

MACRO NOR2_Z3
    CLASS CORE ;
    FOREIGN NOR2_Z3 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.420 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.565 0.150 1.89 0.54 ;
        RECT 1.395 0.150 1.98 0.28 ;
        RECT 1.565 0.505 2.67 0.57 ;
        RECT 2.410 0.505 2.735 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.710 0.340 1.295 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.150 0.340 2.735 0.405 ;
        END
    END b
END NOR2_Z3

MACRO NOR2_Z4
    CLASS CORE ;
    FOREIGN NOR2_Z4 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.740 0.150 2.065 0.54 ;
        RECT 1.550 0.150 2.2 0.28 ;
        RECT 1.740 0.505 2.975 0.57 ;
        RECT 2.675 0.505 3.0 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.790 0.340 1.44 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.390 0.340 3.04 0.405 ;
        END
    END b
END NOR2_Z4

MACRO NOR2_Z6
    CLASS CORE ;
    FOREIGN NOR2_Z6 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.085 0.150 2.475 0.54 ;
        RECT 1.860 0.150 2.64 0.28 ;
        RECT 2.085 0.505 3.58 0.57 ;
        RECT 3.210 0.505 3.6 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.945 0.340 1.725 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.865 0.340 3.645 0.405 ;
        END
    END b
END NOR2_Z6

MACRO NOR2_Z8
    CLASS CORE ;
    FOREIGN NOR2_Z8 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.940 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.260 0.150 2.715 0.54 ;
        RECT 2.015 0.150 2.86 0.28 ;
        RECT 2.260 0.505 3.885 0.57 ;
        RECT 3.480 0.505 3.935 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.025 0.340 1.87 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.105 0.340 3.95 0.405 ;
        END
    END b
END NOR2_Z8

MACRO NOR2_Z10
    CLASS CORE ;
    FOREIGN NOR2_Z10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.700 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.605 0.150 3.125 0.54 ;
        RECT 2.325 0.150 3.365 0.28 ;
        RECT 2.605 0.505 4.49 0.57 ;
        RECT 4.015 0.505 4.535 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.180 0.340 2.09 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.580 0.340 4.49 0.405 ;
        END
    END b
END NOR2_Z10

MACRO NOR2_Z20
    CLASS CORE ;
    FOREIGN NOR2_Z20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.475 0.150 4.125 0.54 ;
        RECT 3.100 0.150 4.465 0.28 ;
        RECT 3.475 0.505 6.01 0.57 ;
        RECT 5.350 0.505 6.0 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.575 0.340 2.81 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.775 0.340 6.01 0.405 ;
        END
    END b
END NOR2_Z20

MACRO NOR2_Z40
    CLASS CORE ;
    FOREIGN NOR2_Z40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.865 0.150 5.775 0.54 ;
        RECT 4.340 0.150 6.225 0.28 ;
        RECT 4.865 0.505 8.375 0.57 ;
        RECT 7.490 0.505 8.4 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.205 0.340 3.96 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.685 0.340 8.44 0.405 ;
        END
    END b
END NOR2_Z40

MACRO NOR2_Z80
    CLASS CORE ;
    FOREIGN NOR2_Z80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.440 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.605 0.150 7.84 0.54 ;
        RECT 5.890 0.150 8.425 0.28 ;
        RECT 6.605 0.505 11.415 0.57 ;
        RECT 10.165 0.505 11.4 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.995 0.340 5.4 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 9.075 0.340 11.48 0.405 ;
        END
    END b
END NOR2_Z80

MACRO NOR3_X1
    CLASS CORE ;
    FOREIGN NOR3_X1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.140 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.420 0.130 0.485 0.39 ;
        RECT 0.420 0.340 0.94 0.405 ;
        RECT 0.870 0.130 0.935 1.625 ;
        RECT 0.870 0.545 0.935 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.085 0.365 0.28 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.415 0.430 0.545 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.645 0.430 0.775 0.56 ;
        END
    END c
END NOR3_X1

MACRO NOR3_X2
    CLASS CORE ;
    FOREIGN NOR3_X2 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.980 0.130 1.175 0.39 ;
        RECT 0.980 0.340 2.215 0.405 ;
        RECT 2.030 0.130 2.225 1.625 ;
        RECT 2.030 0.545 2.225 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.195 0.365 0.65 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.975 0.430 1.3 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.505 0.430 1.83 0.56 ;
        END
    END c
END NOR3_X2

MACRO NOR3_X3
    CLASS CORE ;
    FOREIGN NOR3_X3 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.420 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.260 0.130 1.52 0.39 ;
        RECT 1.260 0.340 2.82 0.405 ;
        RECT 2.610 0.130 2.87 1.625 ;
        RECT 2.610 0.545 2.87 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.250 0.365 0.77 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.250 0.430 1.705 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.935 0.430 2.39 0.56 ;
        END
    END c
END NOR3_X3

MACRO NOR3_X4
    CLASS CORE ;
    FOREIGN NOR3_X4 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.400 0.130 1.66 0.39 ;
        RECT 1.400 0.340 3.155 0.405 ;
        RECT 2.900 0.130 3.16 1.625 ;
        RECT 2.900 0.545 3.16 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.280 0.365 0.865 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.430 1.845 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.150 0.430 2.67 0.56 ;
        END
    END c
END NOR3_X4

MACRO NOR3_X6
    CLASS CORE ;
    FOREIGN NOR3_X6 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.680 0.130 2.005 0.39 ;
        RECT 1.680 0.340 3.76 0.405 ;
        RECT 3.480 0.130 3.805 1.625 ;
        RECT 3.480 0.545 3.805 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.335 0.365 1.05 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.670 0.430 2.255 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.580 0.430 3.165 0.56 ;
        END
    END c
END NOR3_X6

MACRO NOR3_X8
    CLASS CORE ;
    FOREIGN NOR3_X8 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.940 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.820 0.130 2.145 0.39 ;
        RECT 1.820 0.340 4.095 0.405 ;
        RECT 3.770 0.130 4.095 1.625 ;
        RECT 3.770 0.545 4.095 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.365 0.365 1.145 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.805 0.430 2.39 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.795 0.430 3.445 0.56 ;
        END
    END c
END NOR3_X8

MACRO NOR3_X10
    CLASS CORE ;
    FOREIGN NOR3_X10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.700 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.100 0.130 2.49 0.39 ;
        RECT 2.100 0.340 4.765 0.405 ;
        RECT 4.350 0.130 4.74 1.625 ;
        RECT 4.350 0.545 4.74 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.420 0.365 1.33 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.085 0.430 2.8 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.225 0.430 3.94 0.56 ;
        END
    END c
END NOR3_X10

MACRO NOR3_X20
    CLASS CORE ;
    FOREIGN NOR3_X20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.800 0.130 3.32 0.39 ;
        RECT 2.800 0.340 6.31 0.405 ;
        RECT 5.800 0.130 6.32 1.625 ;
        RECT 5.800 0.545 6.32 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.560 0.365 1.795 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.780 0.430 3.69 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.300 0.430 5.275 0.56 ;
        END
    END c
END NOR3_X20

MACRO NOR3_X40
    CLASS CORE ;
    FOREIGN NOR3_X40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.920 0.130 4.635 0.39 ;
        RECT 3.920 0.340 8.86 0.405 ;
        RECT 8.120 0.130 8.835 1.625 ;
        RECT 8.120 0.545 8.9 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.785 0.365 2.475 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.890 0.430 5.19 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.020 0.430 7.385 0.56 ;
        END
    END c
END NOR3_X40

MACRO NOR3_X80
    CLASS CORE ;
    FOREIGN NOR3_X80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.440 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.320 0.130 6.295 0.39 ;
        RECT 5.320 0.340 12.015 0.405 ;
        RECT 11.020 0.130 11.995 1.625 ;
        RECT 11.020 0.545 12.06 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.065 0.365 3.405 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.280 0.430 7.035 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.170 0.430 10.055 0.56 ;
        END
    END c
END NOR3_X80

MACRO NOR3_Y1
    CLASS CORE ;
    FOREIGN NOR3_Y1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.140 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.420 0.130 0.485 0.39 ;
        RECT 0.420 0.340 0.94 0.405 ;
        RECT 0.870 0.130 0.935 1.625 ;
        RECT 0.870 0.545 0.935 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.085 0.365 0.28 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.415 0.430 0.545 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.645 0.430 0.775 0.56 ;
        END
    END c
END NOR3_Y1

MACRO NOR3_Y2
    CLASS CORE ;
    FOREIGN NOR3_Y2 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.980 0.130 1.175 0.39 ;
        RECT 0.980 0.340 2.215 0.405 ;
        RECT 2.030 0.130 2.225 1.625 ;
        RECT 2.030 0.545 2.225 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.195 0.365 0.65 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.975 0.430 1.3 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.505 0.430 1.83 0.56 ;
        END
    END c
END NOR3_Y2

MACRO NOR3_Y3
    CLASS CORE ;
    FOREIGN NOR3_Y3 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.420 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.260 0.130 1.52 0.39 ;
        RECT 1.260 0.340 2.82 0.405 ;
        RECT 2.610 0.130 2.87 1.625 ;
        RECT 2.610 0.545 2.87 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.250 0.365 0.77 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.250 0.430 1.705 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.935 0.430 2.39 0.56 ;
        END
    END c
END NOR3_Y3

MACRO NOR3_Y4
    CLASS CORE ;
    FOREIGN NOR3_Y4 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.400 0.130 1.66 0.39 ;
        RECT 1.400 0.340 3.155 0.405 ;
        RECT 2.900 0.130 3.16 1.625 ;
        RECT 2.900 0.545 3.16 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.280 0.365 0.865 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.430 1.845 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.150 0.430 2.67 0.56 ;
        END
    END c
END NOR3_Y4

MACRO NOR3_Y6
    CLASS CORE ;
    FOREIGN NOR3_Y6 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.680 0.130 2.005 0.39 ;
        RECT 1.680 0.340 3.76 0.405 ;
        RECT 3.480 0.130 3.805 1.625 ;
        RECT 3.480 0.545 3.805 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.335 0.365 1.05 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.670 0.430 2.255 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.580 0.430 3.165 0.56 ;
        END
    END c
END NOR3_Y6

MACRO NOR3_Y8
    CLASS CORE ;
    FOREIGN NOR3_Y8 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.940 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.820 0.130 2.145 0.39 ;
        RECT 1.820 0.340 4.095 0.405 ;
        RECT 3.770 0.130 4.095 1.625 ;
        RECT 3.770 0.545 4.095 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.365 0.365 1.145 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.805 0.430 2.39 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.795 0.430 3.445 0.56 ;
        END
    END c
END NOR3_Y8

MACRO NOR3_Y10
    CLASS CORE ;
    FOREIGN NOR3_Y10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.700 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.100 0.130 2.49 0.39 ;
        RECT 2.100 0.340 4.765 0.405 ;
        RECT 4.350 0.130 4.74 1.625 ;
        RECT 4.350 0.545 4.74 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.420 0.365 1.33 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.085 0.430 2.8 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.225 0.430 3.94 0.56 ;
        END
    END c
END NOR3_Y10

MACRO NOR3_Y20
    CLASS CORE ;
    FOREIGN NOR3_Y20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.800 0.130 3.32 0.39 ;
        RECT 2.800 0.340 6.31 0.405 ;
        RECT 5.800 0.130 6.32 1.625 ;
        RECT 5.800 0.545 6.32 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.560 0.365 1.795 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.780 0.430 3.69 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.300 0.430 5.275 0.56 ;
        END
    END c
END NOR3_Y20

MACRO NOR3_Y40
    CLASS CORE ;
    FOREIGN NOR3_Y40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.920 0.130 4.635 0.39 ;
        RECT 3.920 0.340 8.86 0.405 ;
        RECT 8.120 0.130 8.835 1.625 ;
        RECT 8.120 0.545 8.9 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.785 0.365 2.475 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.890 0.430 5.19 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.020 0.430 7.385 0.56 ;
        END
    END c
END NOR3_Y40

MACRO NOR3_Y80
    CLASS CORE ;
    FOREIGN NOR3_Y80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.440 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.320 0.130 6.295 0.39 ;
        RECT 5.320 0.340 12.015 0.405 ;
        RECT 11.020 0.130 11.995 1.625 ;
        RECT 11.020 0.545 12.06 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.065 0.365 3.405 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.280 0.430 7.035 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.170 0.430 10.055 0.56 ;
        END
    END c
END NOR3_Y80

MACRO NOR3_Z1
    CLASS CORE ;
    FOREIGN NOR3_Z1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.140 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.420 0.130 0.485 0.39 ;
        RECT 0.420 0.340 0.94 0.405 ;
        RECT 0.870 0.130 0.935 1.625 ;
        RECT 0.870 0.545 0.935 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.085 0.365 0.28 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.415 0.430 0.545 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.645 0.430 0.775 0.56 ;
        END
    END c
END NOR3_Z1

MACRO NOR3_Z2
    CLASS CORE ;
    FOREIGN NOR3_Z2 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.980 0.130 1.175 0.39 ;
        RECT 0.980 0.340 2.215 0.405 ;
        RECT 2.030 0.130 2.225 1.625 ;
        RECT 2.030 0.545 2.225 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.195 0.365 0.65 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.975 0.430 1.3 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.505 0.430 1.83 0.56 ;
        END
    END c
END NOR3_Z2

MACRO NOR3_Z3
    CLASS CORE ;
    FOREIGN NOR3_Z3 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.420 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.260 0.130 1.52 0.39 ;
        RECT 1.260 0.340 2.82 0.405 ;
        RECT 2.610 0.130 2.87 1.625 ;
        RECT 2.610 0.545 2.87 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.250 0.365 0.77 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.250 0.430 1.705 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.935 0.430 2.39 0.56 ;
        END
    END c
END NOR3_Z3

MACRO NOR3_Z4
    CLASS CORE ;
    FOREIGN NOR3_Z4 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.400 0.130 1.66 0.39 ;
        RECT 1.400 0.340 3.155 0.405 ;
        RECT 2.900 0.130 3.16 1.625 ;
        RECT 2.900 0.545 3.16 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.280 0.365 0.865 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.430 1.845 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.150 0.430 2.67 0.56 ;
        END
    END c
END NOR3_Z4

MACRO NOR3_Z6
    CLASS CORE ;
    FOREIGN NOR3_Z6 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.680 0.130 2.005 0.39 ;
        RECT 1.680 0.340 3.76 0.405 ;
        RECT 3.480 0.130 3.805 1.625 ;
        RECT 3.480 0.545 3.805 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.335 0.365 1.05 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.670 0.430 2.255 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.580 0.430 3.165 0.56 ;
        END
    END c
END NOR3_Z6

MACRO NOR3_Z8
    CLASS CORE ;
    FOREIGN NOR3_Z8 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.940 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.820 0.130 2.145 0.39 ;
        RECT 1.820 0.340 4.095 0.405 ;
        RECT 3.770 0.130 4.095 1.625 ;
        RECT 3.770 0.545 4.095 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.365 0.365 1.145 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.805 0.430 2.39 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.795 0.430 3.445 0.56 ;
        END
    END c
END NOR3_Z8

MACRO NOR3_Z10
    CLASS CORE ;
    FOREIGN NOR3_Z10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.700 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.100 0.130 2.49 0.39 ;
        RECT 2.100 0.340 4.765 0.405 ;
        RECT 4.350 0.130 4.74 1.625 ;
        RECT 4.350 0.545 4.74 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.420 0.365 1.33 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.085 0.430 2.8 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.225 0.430 3.94 0.56 ;
        END
    END c
END NOR3_Z10

MACRO NOR3_Z20
    CLASS CORE ;
    FOREIGN NOR3_Z20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.800 0.130 3.32 0.39 ;
        RECT 2.800 0.340 6.31 0.405 ;
        RECT 5.800 0.130 6.32 1.625 ;
        RECT 5.800 0.545 6.32 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.560 0.365 1.795 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.780 0.430 3.69 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.300 0.430 5.275 0.56 ;
        END
    END c
END NOR3_Z20

MACRO NOR3_Z40
    CLASS CORE ;
    FOREIGN NOR3_Z40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.920 0.130 4.635 0.39 ;
        RECT 3.920 0.340 8.86 0.405 ;
        RECT 8.120 0.130 8.835 1.625 ;
        RECT 8.120 0.545 8.9 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.785 0.365 2.475 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.890 0.430 5.19 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.020 0.430 7.385 0.56 ;
        END
    END c
END NOR3_Z40

MACRO NOR3_Z80
    CLASS CORE ;
    FOREIGN NOR3_Z80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.440 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.320 0.130 6.295 0.39 ;
        RECT 5.320 0.340 12.015 0.405 ;
        RECT 11.020 0.130 11.995 1.625 ;
        RECT 11.020 0.545 12.06 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.065 0.365 3.405 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.280 0.430 7.035 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.170 0.430 10.055 0.56 ;
        END
    END c
END NOR3_Z80

MACRO NOR4_X1
    CLASS CORE ;
    FOREIGN NOR4_X1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.520 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.465 0.090 0.53 1.455 ;
        RECT 0.465 0.090 0.79 0.155 ;
        RECT 0.715 0.090 0.78 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.145 0.530 1.34 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.890 0.530 1.085 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.045 0.530 0.305 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.635 0.530 0.83 0.66 ;
        END
    END d
END NOR4_X1

MACRO NOR4_X2
    CLASS CORE ;
    FOREIGN NOR4_X2 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.040 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.925 0.090 1.12 1.455 ;
        RECT 0.925 0.090 1.575 0.155 ;
        RECT 1.425 0.090 1.62 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.285 0.530 2.61 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.780 0.530 2.105 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.085 0.530 0.605 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.275 0.530 1.6 0.66 ;
        END
    END d
END NOR4_X2

MACRO NOR4_X3
    CLASS CORE ;
    FOREIGN NOR4_X3 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.160 0.090 1.355 1.455 ;
        RECT 1.160 0.090 2.005 0.155 ;
        RECT 1.785 0.090 1.98 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.860 0.530 3.25 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.225 0.530 2.615 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.110 0.530 0.76 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.590 0.530 1.98 0.66 ;
        END
    END d
END NOR4_X3

MACRO NOR4_X4
    CLASS CORE ;
    FOREIGN NOR4_X4 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.090 1.65 1.455 ;
        RECT 1.390 0.090 2.43 0.155 ;
        RECT 2.140 0.090 2.4 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.430 0.530 3.95 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.670 0.530 3.19 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.130 0.530 0.91 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.910 0.530 2.43 0.66 ;
        END
    END d
END NOR4_X4

MACRO NOR4_X6
    CLASS CORE ;
    FOREIGN NOR4_X6 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.620 0.090 1.945 1.455 ;
        RECT 1.620 0.090 2.79 0.155 ;
        RECT 2.495 0.090 2.82 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.000 0.530 4.585 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.115 0.530 3.7 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.150 0.530 1.06 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.230 0.530 2.815 0.66 ;
        END
    END d
END NOR4_X6

MACRO NOR4_X8
    CLASS CORE ;
    FOREIGN NOR4_X8 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.080 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.855 0.090 2.18 1.455 ;
        RECT 1.855 0.090 3.22 0.155 ;
        RECT 2.855 0.090 3.18 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.575 0.530 5.225 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.560 0.530 4.21 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.175 0.530 1.215 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.545 0.530 3.195 0.66 ;
        END
    END d
END NOR4_X8

MACRO NOR4_X10
    CLASS CORE ;
    FOREIGN NOR4_X10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.460 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.970 0.090 2.36 1.455 ;
        RECT 1.970 0.090 3.4 0.155 ;
        RECT 3.030 0.090 3.42 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.860 0.530 5.575 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.785 0.530 4.5 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.185 0.530 1.29 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.705 0.530 3.42 0.66 ;
        END
    END d
END NOR4_X10

MACRO NOR4_X20
    CLASS CORE ;
    FOREIGN NOR4_X20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.740 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.665 0.090 3.185 1.455 ;
        RECT 2.665 0.090 4.615 0.155 ;
        RECT 4.100 0.090 4.62 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.575 0.530 7.55 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.115 0.530 6.09 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.250 0.530 1.68 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.660 0.530 4.635 0.66 ;
        END
    END d
END NOR4_X20

MACRO NOR4_X40
    CLASS CORE ;
    FOREIGN NOR4_X40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.780 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.590 0.090 4.24 1.455 ;
        RECT 3.590 0.090 6.19 0.155 ;
        RECT 5.530 0.090 6.18 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.860 0.530 10.16 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.895 0.530 8.195 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.335 0.530 2.285 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.935 0.530 6.235 0.66 ;
        END
    END d
END NOR4_X40

MACRO NOR4_X80
    CLASS CORE ;
    FOREIGN NOR4_X80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.340 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.980 0.090 5.89 1.455 ;
        RECT 4.980 0.090 8.62 0.155 ;
        RECT 7.670 0.090 8.58 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 12.290 0.530 14.11 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 9.565 0.530 11.385 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.465 0.530 3.195 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.845 0.530 8.665 0.66 ;
        END
    END d
END NOR4_X80

MACRO NOR4_Y1
    CLASS CORE ;
    FOREIGN NOR4_Y1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.520 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.465 0.090 0.53 1.455 ;
        RECT 0.465 0.090 0.79 0.155 ;
        RECT 0.715 0.090 0.78 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.145 0.530 1.34 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.890 0.530 1.085 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.045 0.530 0.305 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.635 0.530 0.83 0.66 ;
        END
    END d
END NOR4_Y1

MACRO NOR4_Y2
    CLASS CORE ;
    FOREIGN NOR4_Y2 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.040 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.925 0.090 1.12 1.455 ;
        RECT 0.925 0.090 1.575 0.155 ;
        RECT 1.425 0.090 1.62 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.285 0.530 2.61 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.780 0.530 2.105 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.085 0.530 0.605 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.275 0.530 1.6 0.66 ;
        END
    END d
END NOR4_Y2

MACRO NOR4_Y3
    CLASS CORE ;
    FOREIGN NOR4_Y3 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.160 0.090 1.355 1.455 ;
        RECT 1.160 0.090 2.005 0.155 ;
        RECT 1.785 0.090 1.98 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.860 0.530 3.25 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.225 0.530 2.615 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.110 0.530 0.76 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.590 0.530 1.98 0.66 ;
        END
    END d
END NOR4_Y3

MACRO NOR4_Y4
    CLASS CORE ;
    FOREIGN NOR4_Y4 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.090 1.65 1.455 ;
        RECT 1.390 0.090 2.43 0.155 ;
        RECT 2.140 0.090 2.4 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.430 0.530 3.95 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.670 0.530 3.19 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.130 0.530 0.91 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.910 0.530 2.43 0.66 ;
        END
    END d
END NOR4_Y4

MACRO NOR4_Y6
    CLASS CORE ;
    FOREIGN NOR4_Y6 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.620 0.090 1.945 1.455 ;
        RECT 1.620 0.090 2.79 0.155 ;
        RECT 2.495 0.090 2.82 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.000 0.530 4.585 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.115 0.530 3.7 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.150 0.530 1.06 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.230 0.530 2.815 0.66 ;
        END
    END d
END NOR4_Y6

MACRO NOR4_Y8
    CLASS CORE ;
    FOREIGN NOR4_Y8 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.080 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.855 0.090 2.18 1.455 ;
        RECT 1.855 0.090 3.22 0.155 ;
        RECT 2.855 0.090 3.18 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.575 0.530 5.225 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.560 0.530 4.21 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.175 0.530 1.215 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.545 0.530 3.195 0.66 ;
        END
    END d
END NOR4_Y8

MACRO NOR4_Y10
    CLASS CORE ;
    FOREIGN NOR4_Y10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.460 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.970 0.090 2.36 1.455 ;
        RECT 1.970 0.090 3.4 0.155 ;
        RECT 3.030 0.090 3.42 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.860 0.530 5.575 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.785 0.530 4.5 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.185 0.530 1.29 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.705 0.530 3.42 0.66 ;
        END
    END d
END NOR4_Y10

MACRO NOR4_Y20
    CLASS CORE ;
    FOREIGN NOR4_Y20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.740 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.665 0.090 3.185 1.455 ;
        RECT 2.665 0.090 4.615 0.155 ;
        RECT 4.100 0.090 4.62 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.575 0.530 7.55 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.115 0.530 6.09 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.250 0.530 1.68 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.660 0.530 4.635 0.66 ;
        END
    END d
END NOR4_Y20

MACRO NOR4_Y40
    CLASS CORE ;
    FOREIGN NOR4_Y40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.780 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.590 0.090 4.24 1.455 ;
        RECT 3.590 0.090 6.19 0.155 ;
        RECT 5.530 0.090 6.18 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.860 0.530 10.16 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.895 0.530 8.195 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.335 0.530 2.285 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.935 0.530 6.235 0.66 ;
        END
    END d
END NOR4_Y40

MACRO NOR4_Y80
    CLASS CORE ;
    FOREIGN NOR4_Y80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.340 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.980 0.090 5.89 1.455 ;
        RECT 4.980 0.090 8.62 0.155 ;
        RECT 7.670 0.090 8.58 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 12.290 0.530 14.11 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 9.565 0.530 11.385 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.465 0.530 3.195 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.845 0.530 8.665 0.66 ;
        END
    END d
END NOR4_Y80

MACRO NOR4_Z1
    CLASS CORE ;
    FOREIGN NOR4_Z1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.520 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.465 0.090 0.53 1.455 ;
        RECT 0.465 0.090 0.79 0.155 ;
        RECT 0.715 0.090 0.78 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.145 0.530 1.34 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.890 0.530 1.085 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.045 0.530 0.305 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.635 0.530 0.83 0.66 ;
        END
    END d
END NOR4_Z1

MACRO NOR4_Z2
    CLASS CORE ;
    FOREIGN NOR4_Z2 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.040 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.925 0.090 1.12 1.455 ;
        RECT 0.925 0.090 1.575 0.155 ;
        RECT 1.425 0.090 1.62 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.285 0.530 2.61 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.780 0.530 2.105 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.085 0.530 0.605 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.275 0.530 1.6 0.66 ;
        END
    END d
END NOR4_Z2

MACRO NOR4_Z3
    CLASS CORE ;
    FOREIGN NOR4_Z3 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.160 0.090 1.355 1.455 ;
        RECT 1.160 0.090 2.005 0.155 ;
        RECT 1.785 0.090 1.98 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.860 0.530 3.25 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.225 0.530 2.615 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.110 0.530 0.76 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.590 0.530 1.98 0.66 ;
        END
    END d
END NOR4_Z3

MACRO NOR4_Z4
    CLASS CORE ;
    FOREIGN NOR4_Z4 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.090 1.65 1.455 ;
        RECT 1.390 0.090 2.43 0.155 ;
        RECT 2.140 0.090 2.4 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.430 0.530 3.95 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.670 0.530 3.19 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.130 0.530 0.91 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.910 0.530 2.43 0.66 ;
        END
    END d
END NOR4_Z4

MACRO NOR4_Z6
    CLASS CORE ;
    FOREIGN NOR4_Z6 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.620 0.090 1.945 1.455 ;
        RECT 1.620 0.090 2.79 0.155 ;
        RECT 2.495 0.090 2.82 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.000 0.530 4.585 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.115 0.530 3.7 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.150 0.530 1.06 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.230 0.530 2.815 0.66 ;
        END
    END d
END NOR4_Z6

MACRO NOR4_Z8
    CLASS CORE ;
    FOREIGN NOR4_Z8 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.080 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.855 0.090 2.18 1.455 ;
        RECT 1.855 0.090 3.22 0.155 ;
        RECT 2.855 0.090 3.18 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.575 0.530 5.225 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.560 0.530 4.21 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.175 0.530 1.215 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.545 0.530 3.195 0.66 ;
        END
    END d
END NOR4_Z8

MACRO NOR4_Z10
    CLASS CORE ;
    FOREIGN NOR4_Z10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.460 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.970 0.090 2.36 1.455 ;
        RECT 1.970 0.090 3.4 0.155 ;
        RECT 3.030 0.090 3.42 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.860 0.530 5.575 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.785 0.530 4.5 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.185 0.530 1.29 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.705 0.530 3.42 0.66 ;
        END
    END d
END NOR4_Z10

MACRO NOR4_Z20
    CLASS CORE ;
    FOREIGN NOR4_Z20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.740 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.665 0.090 3.185 1.455 ;
        RECT 2.665 0.090 4.615 0.155 ;
        RECT 4.100 0.090 4.62 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.575 0.530 7.55 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.115 0.530 6.09 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.250 0.530 1.68 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.660 0.530 4.635 0.66 ;
        END
    END d
END NOR4_Z20

MACRO NOR4_Z40
    CLASS CORE ;
    FOREIGN NOR4_Z40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.780 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.590 0.090 4.24 1.455 ;
        RECT 3.590 0.090 6.19 0.155 ;
        RECT 5.530 0.090 6.18 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.860 0.530 10.16 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.895 0.530 8.195 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.335 0.530 2.285 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.935 0.530 6.235 0.66 ;
        END
    END d
END NOR4_Z40

MACRO NOR4_Z80
    CLASS CORE ;
    FOREIGN NOR4_Z80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.340 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.980 0.090 5.89 1.455 ;
        RECT 4.980 0.090 8.62 0.155 ;
        RECT 7.670 0.090 8.58 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 12.290 0.530 14.11 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 9.565 0.530 11.385 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.465 0.530 3.195 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.845 0.530 8.665 0.66 ;
        END
    END d
END NOR4_Z80

MACRO DFF_X80
    CLASS CORE ;
    FOREIGN DFF_X80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.500 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.190 0.150 0.45 1.58 ;
        RECT 0.190 0.635 0.775 0.7 ;
        RECT 0.190 1.140 1.62 1.205 ;
        END
    END q
    PIN ck
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.240 0.990 5.5 1.38 ;
        RECT 5.240 0.990 5.565 1.185 ;
        RECT 1.815 0.640 2.075 0.835 ;
        RECT 1.565 0.780 2.02 0.845 ;
        RECT 1.815 0.640 3.505 0.705 ;
        RECT 2.815 0.640 3.53 0.835 ;
        RECT 4.330 0.705 4.785 0.835 ;
        RECT 2.815 0.790 4.83 0.855 ;
        RECT 4.580 0.705 4.84 1.03 ;
        RECT 4.580 1.015 5.685 1.08 ;
        RECT 5.190 1.015 5.645 1.145 ;
        RECT 5.240 1.290 5.5 1.485 ;
        RECT 7.940 0.775 8.46 0.84 ;
        RECT 8.240 0.775 8.5 1.49 ;
        RECT 5.240 1.470 8.49 1.535 ;
        RECT 5.240 1.315 5.5 1.38 ;
        RECT 5.315 1.110 5.575 1.175 ;
        RECT 5.315 1.015 5.575 1.08 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.705 0.720 8.965 0.785 ;
        END
    END d
END DFF_X80

MACRO TIEH_X1
    CLASS CORE ;
    FOREIGN TIEH_X1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.520 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
				USE SIGNAL ;
        PORT
        LAYER metal1 ;
        RECT 0.925 0.150 1.12 1.255 ;
        RECT 0.835 0.150 1.225 0.28 ;
        END
    END o
END TIEH_X1

MACRO block_9x9_0
 CLASS BLOCK ;
 FOREIGN block_9x9_0 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 3.42 BY 1.71 ;
 SYMMETRY X Y ;
 OBS
  LAYER metal1 ;
   RECT 0 0 3.42 1.71 ;
  LAYER via1 ;
   RECT 0 0 3.42 1.71 ;
  LAYER metal2 ;
   RECT 0 0 3.42 1.71 ;
  LAYER via2 ;
   RECT 0 0 3.42 1.71 ;
  LAYER metal3 ;
   RECT 0 0 3.42 1.71 ;
  LAYER via3 ;
   RECT 0 0 3.42 1.71 ;
  LAYER metal4 ;
   RECT 0 0 3.42 1.71 ;
 END
END block_9x9_0

MACRO block_414x2007_358
 CLASS BLOCK ;
 FOREIGN block_414x2007_358 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 157.32 BY 381.33 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 371.355 26.885 371.925 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 367.175 26.885 367.745 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 346.845 26.885 347.415 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 342.665 26.885 343.235 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 322.335 26.885 322.905 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 318.155 26.885 318.725 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 279.585 26.885 280.155 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 275.405 26.885 275.975 ;
  END
 END o7
 PIN o8
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 255.075 26.885 255.645 ;
  END
 END o8
 PIN o9
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 250.895 26.885 251.465 ;
  END
 END o9
 PIN o10
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 230.565 26.885 231.135 ;
  END
 END o10
 PIN o11
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 226.385 26.885 226.955 ;
  END
 END o11
 PIN o12
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 206.055 26.885 206.625 ;
  END
 END o12
 PIN o13
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 177.745 26.885 178.315 ;
  END
 END o13
 PIN o14
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 157.415 26.885 157.985 ;
  END
 END o14
 PIN o15
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 153.235 26.885 153.805 ;
  END
 END o15
 PIN o16
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 246.905 26.885 247.475 ;
  END
 END o16
 PIN o17
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 173.755 26.885 174.325 ;
  END
 END o17
 PIN o18
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 338.675 26.885 339.245 ;
  END
 END o18
 PIN o19
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 314.165 26.885 314.735 ;
  END
 END o19
 PIN o20
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 149.245 26.885 149.815 ;
  END
 END o20
 PIN o21
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 271.415 26.885 271.985 ;
  END
 END o21
 PIN o22
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 222.395 26.885 222.965 ;
  END
 END o22
 PIN o23
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 363.185 26.885 363.755 ;
  END
 END o23
 PIN o24
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 77.805 26.885 78.375 ;
  END
 END o24
 PIN o25
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 124.735 26.885 125.305 ;
  END
 END o25
 PIN o26
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 301.815 26.885 302.385 ;
  END
 END o26
 PIN o27
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 259.065 26.885 259.635 ;
  END
 END o27
 PIN o28
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 145.065 26.885 145.635 ;
  END
 END o28
 PIN o29
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 112.385 26.885 112.955 ;
  END
 END o29
 PIN o30
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 132.905 26.885 133.475 ;
  END
 END o30
 PIN o31
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 81.985 26.885 82.555 ;
  END
 END o31
 PIN o32
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 334.495 26.885 335.065 ;
  END
 END o32
 PIN o33
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 165.585 26.885 166.155 ;
  END
 END o33
 PIN o34
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 161.405 26.885 161.975 ;
  END
 END o34
 PIN o35
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 169.575 26.885 170.145 ;
  END
 END o35
 PIN o36
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 73.815 26.885 74.385 ;
  END
 END o36
 PIN o37
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 69.635 26.885 70.205 ;
  END
 END o37
 PIN o38
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 65.645 26.885 66.215 ;
  END
 END o38
 PIN o39
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 8.455 26.885 9.025 ;
  END
 END o39
 PIN o40
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 12.445 26.885 13.015 ;
  END
 END o40
 PIN o41
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 45.125 26.885 45.695 ;
  END
 END o41
 PIN o42
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 49.305 26.885 49.875 ;
  END
 END o42
 PIN o43
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 36.955 26.885 37.525 ;
  END
 END o43
 PIN o44
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 41.135 26.885 41.705 ;
  END
 END o44
 PIN o45
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 116.565 26.885 117.135 ;
  END
 END o45
 PIN o46
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 359.005 26.885 359.575 ;
  END
 END o46
 PIN o47
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 350.835 26.885 351.405 ;
  END
 END o47
 PIN o48
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 326.325 26.885 326.895 ;
  END
 END o48
 PIN o49
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 263.245 26.885 263.815 ;
  END
 END o49
 PIN o50
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 24.795 26.885 25.365 ;
  END
 END o50
 PIN o51
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 53.295 26.885 53.865 ;
  END
 END o51
 PIN o52
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 234.555 26.885 235.125 ;
  END
 END o52
 PIN o53
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 4.275 26.885 4.845 ;
  END
 END o53
 PIN o54
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 128.725 26.885 129.295 ;
  END
 END o54
 PIN o55
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 214.225 26.885 214.795 ;
  END
 END o55
 PIN o56
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 32.965 26.885 33.535 ;
  END
 END o56
 PIN o57
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 57.475 26.885 58.045 ;
  END
 END o57
 PIN o58
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 28.785 26.885 29.355 ;
  END
 END o58
 PIN o59
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 104.215 26.885 104.785 ;
  END
 END o59
 PIN o60
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 61.465 26.885 62.035 ;
  END
 END o60
 PIN o61
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 120.555 26.885 121.125 ;
  END
 END o61
 PIN o62
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 242.725 26.885 243.295 ;
  END
 END o62
 PIN o63
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 238.735 26.885 239.305 ;
  END
 END o63
 PIN o64
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 355.015 26.885 355.585 ;
  END
 END o64
 PIN o65
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 108.395 26.885 108.965 ;
  END
 END o65
 PIN o66
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 141.075 26.885 141.645 ;
  END
 END o66
 PIN o67
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 136.895 26.885 137.465 ;
  END
 END o67
 PIN o68
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 218.215 26.885 218.785 ;
  END
 END o68
 PIN o69
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 267.235 26.885 267.805 ;
  END
 END o69
 PIN o70
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 305.995 26.885 306.565 ;
  END
 END o70
 PIN o71
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 309.985 26.885 310.555 ;
  END
 END o71
 PIN o72
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 330.505 26.885 331.075 ;
  END
 END o72
 PIN o73
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 20.615 26.885 21.185 ;
  END
 END o73
 PIN o74
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 16.625 26.885 17.195 ;
  END
 END o74
 PIN o75
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 210.045 26.885 210.615 ;
  END
 END o75
 PIN o76
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 375.345 26.885 375.915 ;
  END
 END o76
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 180.785 3.705 181.355 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 197.885 3.705 198.455 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 186.105 3.705 186.675 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 181.165 4.465 181.735 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 180.405 4.465 180.975 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 180.025 3.705 180.595 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 189.715 3.705 190.285 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 202.825 3.705 203.395 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 197.125 3.705 197.695 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 199.215 3.705 199.785 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 201.685 3.705 202.255 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 203.205 4.465 203.775 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 13.015 179.645 13.585 180.215 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 13.015 192.945 13.585 193.515 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 2.565 26.885 3.135 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 6.745 26.885 7.315 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 43.415 26.885 43.985 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 47.595 26.885 48.165 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 51.585 26.885 52.155 ;
  END
 END i18
 PIN i19
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 55.765 26.885 56.335 ;
  END
 END i19
 PIN i20
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 59.755 26.885 60.325 ;
  END
 END i20
 PIN i21
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 63.935 26.885 64.505 ;
  END
 END i21
 PIN i22
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 67.925 26.885 68.495 ;
  END
 END i22
 PIN i23
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 72.105 26.885 72.675 ;
  END
 END i23
 PIN i24
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 76.095 26.885 76.665 ;
  END
 END i24
 PIN i25
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 80.275 26.885 80.845 ;
  END
 END i25
 PIN i26
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 10.735 26.885 11.305 ;
  END
 END i26
 PIN i27
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 102.505 26.885 103.075 ;
  END
 END i27
 PIN i28
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 106.685 26.885 107.255 ;
  END
 END i28
 PIN i29
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 110.675 26.885 111.245 ;
  END
 END i29
 PIN i30
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 114.855 26.885 115.425 ;
  END
 END i30
 PIN i31
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 118.845 26.885 119.415 ;
  END
 END i31
 PIN i32
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 123.025 26.885 123.595 ;
  END
 END i32
 PIN i33
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 127.015 26.885 127.585 ;
  END
 END i33
 PIN i34
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 131.195 26.885 131.765 ;
  END
 END i34
 PIN i35
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 135.185 26.885 135.755 ;
  END
 END i35
 PIN i36
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 139.365 26.885 139.935 ;
  END
 END i36
 PIN i37
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 14.915 26.885 15.485 ;
  END
 END i37
 PIN i38
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 143.355 26.885 143.925 ;
  END
 END i38
 PIN i39
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 147.535 26.885 148.105 ;
  END
 END i39
 PIN i40
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 151.525 26.885 152.095 ;
  END
 END i40
 PIN i41
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 155.705 26.885 156.275 ;
  END
 END i41
 PIN i42
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 159.695 26.885 160.265 ;
  END
 END i42
 PIN i43
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 163.875 26.885 164.445 ;
  END
 END i43
 PIN i44
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 167.865 26.885 168.435 ;
  END
 END i44
 PIN i45
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 172.045 26.885 172.615 ;
  END
 END i45
 PIN i46
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 176.035 26.885 176.605 ;
  END
 END i46
 PIN i47
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 207.765 26.885 208.335 ;
  END
 END i47
 PIN i48
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 18.905 26.885 19.475 ;
  END
 END i48
 PIN i49
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 211.755 26.885 212.325 ;
  END
 END i49
 PIN i50
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 215.935 26.885 216.505 ;
  END
 END i50
 PIN i51
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 219.925 26.885 220.495 ;
  END
 END i51
 PIN i52
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 224.105 26.885 224.675 ;
  END
 END i52
 PIN i53
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 228.095 26.885 228.665 ;
  END
 END i53
 PIN i54
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 232.275 26.885 232.845 ;
  END
 END i54
 PIN i55
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 236.265 26.885 236.835 ;
  END
 END i55
 PIN i56
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 240.445 26.885 241.015 ;
  END
 END i56
 PIN i57
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 244.435 26.885 245.005 ;
  END
 END i57
 PIN i58
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 248.615 26.885 249.185 ;
  END
 END i58
 PIN i59
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 23.085 26.885 23.655 ;
  END
 END i59
 PIN i60
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 252.605 26.885 253.175 ;
  END
 END i60
 PIN i61
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 256.785 26.885 257.355 ;
  END
 END i61
 PIN i62
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 260.775 26.885 261.345 ;
  END
 END i62
 PIN i63
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 264.955 26.885 265.525 ;
  END
 END i63
 PIN i64
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 268.945 26.885 269.515 ;
  END
 END i64
 PIN i65
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 273.125 26.885 273.695 ;
  END
 END i65
 PIN i66
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 277.115 26.885 277.685 ;
  END
 END i66
 PIN i67
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 281.295 26.885 281.865 ;
  END
 END i67
 PIN i68
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 303.525 26.885 304.095 ;
  END
 END i68
 PIN i69
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 307.705 26.885 308.275 ;
  END
 END i69
 PIN i70
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 27.075 26.885 27.645 ;
  END
 END i70
 PIN i71
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 311.695 26.885 312.265 ;
  END
 END i71
 PIN i72
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 315.875 26.885 316.445 ;
  END
 END i72
 PIN i73
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 319.865 26.885 320.435 ;
  END
 END i73
 PIN i74
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 324.045 26.885 324.615 ;
  END
 END i74
 PIN i75
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 328.035 26.885 328.605 ;
  END
 END i75
 PIN i76
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 332.215 26.885 332.785 ;
  END
 END i76
 PIN i77
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 336.205 26.885 336.775 ;
  END
 END i77
 PIN i78
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 340.385 26.885 340.955 ;
  END
 END i78
 PIN i79
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 344.375 26.885 344.945 ;
  END
 END i79
 PIN i80
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 348.555 26.885 349.125 ;
  END
 END i80
 PIN i81
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 31.255 26.885 31.825 ;
  END
 END i81
 PIN i82
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 352.545 26.885 353.115 ;
  END
 END i82
 PIN i83
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 356.725 26.885 357.295 ;
  END
 END i83
 PIN i84
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 360.715 26.885 361.285 ;
  END
 END i84
 PIN i85
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 364.895 26.885 365.465 ;
  END
 END i85
 PIN i86
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 368.885 26.885 369.455 ;
  END
 END i86
 PIN i87
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 373.065 26.885 373.635 ;
  END
 END i87
 PIN i88
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 377.055 26.885 377.625 ;
  END
 END i88
 PIN i89
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 35.245 26.885 35.815 ;
  END
 END i89
 PIN i90
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 39.425 26.885 39.995 ;
  END
 END i90
 PIN i91
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 58.045 27.645 58.615 ;
  END
 END i91
 PIN i92
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 62.035 27.645 62.605 ;
  END
 END i92
 PIN i93
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 66.215 27.645 66.785 ;
  END
 END i93
 PIN i94
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 45.695 27.645 46.265 ;
  END
 END i94
 PIN i95
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 49.875 27.645 50.445 ;
  END
 END i95
 PIN i96
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 125.305 27.645 125.875 ;
  END
 END i96
 PIN i97
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 129.295 27.645 129.865 ;
  END
 END i97
 PIN i98
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 133.475 27.645 134.045 ;
  END
 END i98
 PIN i99
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 137.465 27.645 138.035 ;
  END
 END i99
 PIN i100
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 141.645 27.645 142.215 ;
  END
 END i100
 PIN i101
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 258.495 27.645 259.065 ;
  END
 END i101
 PIN i102
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 254.505 27.645 255.075 ;
  END
 END i102
 PIN i103
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 250.325 27.645 250.895 ;
  END
 END i103
 PIN i104
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 246.335 27.645 246.905 ;
  END
 END i104
 PIN i105
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 242.155 27.645 242.725 ;
  END
 END i105
 PIN i106
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 325.755 27.645 326.325 ;
  END
 END i106
 PIN i107
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 321.765 27.645 322.335 ;
  END
 END i107
 PIN i108
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 317.585 27.645 318.155 ;
  END
 END i108
 PIN i109
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 338.105 27.645 338.675 ;
  END
 END i109
 PIN i110
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 333.925 27.645 334.495 ;
  END
 END i110
 PIN i111
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 53.865 27.645 54.435 ;
  END
 END i111
 PIN i112
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 121.125 27.645 121.695 ;
  END
 END i112
 PIN i113
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 262.675 27.645 263.245 ;
  END
 END i113
 PIN i114
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 329.935 27.645 330.505 ;
  END
 END i114
 PIN i115
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 17.955 179.645 18.525 180.215 ;
  END
 END i115
 PIN i116
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 17.955 192.945 18.525 193.515 ;
  END
 END i116
 PIN i117
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 3.135 27.645 3.705 ;
  END
 END i117
 PIN i118
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 7.315 27.645 7.885 ;
  END
 END i118
 PIN i119
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 43.985 27.645 44.555 ;
  END
 END i119
 PIN i120
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 48.165 27.645 48.735 ;
  END
 END i120
 PIN i121
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 52.155 27.645 52.725 ;
  END
 END i121
 PIN i122
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 56.335 27.645 56.905 ;
  END
 END i122
 PIN i123
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 60.325 27.645 60.895 ;
  END
 END i123
 PIN i124
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 64.505 27.645 65.075 ;
  END
 END i124
 PIN i125
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 68.495 27.645 69.065 ;
  END
 END i125
 PIN i126
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 72.675 27.645 73.245 ;
  END
 END i126
 PIN i127
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 76.665 27.645 77.235 ;
  END
 END i127
 PIN i128
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 80.845 27.645 81.415 ;
  END
 END i128
 PIN i129
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 11.305 27.645 11.875 ;
  END
 END i129
 PIN i130
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 103.075 27.645 103.645 ;
  END
 END i130
 PIN i131
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 107.255 27.645 107.825 ;
  END
 END i131
 PIN i132
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 111.245 27.645 111.815 ;
  END
 END i132
 PIN i133
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 115.425 27.645 115.995 ;
  END
 END i133
 PIN i134
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 119.415 27.645 119.985 ;
  END
 END i134
 PIN i135
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 123.595 27.645 124.165 ;
  END
 END i135
 PIN i136
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 127.585 27.645 128.155 ;
  END
 END i136
 PIN i137
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 131.765 27.645 132.335 ;
  END
 END i137
 PIN i138
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 135.755 27.645 136.325 ;
  END
 END i138
 PIN i139
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 139.935 27.645 140.505 ;
  END
 END i139
 PIN i140
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 15.485 27.645 16.055 ;
  END
 END i140
 PIN i141
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 143.925 27.645 144.495 ;
  END
 END i141
 PIN i142
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 148.105 27.645 148.675 ;
  END
 END i142
 PIN i143
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 152.095 27.645 152.665 ;
  END
 END i143
 PIN i144
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 156.275 27.645 156.845 ;
  END
 END i144
 PIN i145
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 160.265 27.645 160.835 ;
  END
 END i145
 PIN i146
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 164.445 27.645 165.015 ;
  END
 END i146
 PIN i147
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 168.435 27.645 169.005 ;
  END
 END i147
 PIN i148
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 172.615 27.645 173.185 ;
  END
 END i148
 PIN i149
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 176.605 27.645 177.175 ;
  END
 END i149
 PIN i150
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 207.195 27.645 207.765 ;
  END
 END i150
 PIN i151
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 19.475 27.645 20.045 ;
  END
 END i151
 PIN i152
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 211.185 27.645 211.755 ;
  END
 END i152
 PIN i153
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 215.365 27.645 215.935 ;
  END
 END i153
 PIN i154
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 219.355 27.645 219.925 ;
  END
 END i154
 PIN i155
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 223.535 27.645 224.105 ;
  END
 END i155
 PIN i156
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 227.525 27.645 228.095 ;
  END
 END i156
 PIN i157
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 231.705 27.645 232.275 ;
  END
 END i157
 PIN i158
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 235.695 27.645 236.265 ;
  END
 END i158
 PIN i159
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 239.875 27.645 240.445 ;
  END
 END i159
 PIN i160
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 243.865 27.645 244.435 ;
  END
 END i160
 PIN i161
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 248.045 27.645 248.615 ;
  END
 END i161
 PIN i162
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 23.655 27.645 24.225 ;
  END
 END i162
 PIN i163
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 252.035 27.645 252.605 ;
  END
 END i163
 PIN i164
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 256.215 27.645 256.785 ;
  END
 END i164
 PIN i165
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 260.205 27.645 260.775 ;
  END
 END i165
 PIN i166
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 264.385 27.645 264.955 ;
  END
 END i166
 PIN i167
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 268.375 27.645 268.945 ;
  END
 END i167
 PIN i168
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 272.555 27.645 273.125 ;
  END
 END i168
 PIN i169
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 276.545 27.645 277.115 ;
  END
 END i169
 PIN i170
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 280.725 27.645 281.295 ;
  END
 END i170
 PIN i171
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 302.955 27.645 303.525 ;
  END
 END i171
 PIN i172
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 307.135 27.645 307.705 ;
  END
 END i172
 PIN i173
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 27.645 27.645 28.215 ;
  END
 END i173
 PIN i174
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 311.125 27.645 311.695 ;
  END
 END i174
 PIN i175
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 315.305 27.645 315.875 ;
  END
 END i175
 PIN i176
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 319.295 27.645 319.865 ;
  END
 END i176
 PIN i177
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 323.475 27.645 324.045 ;
  END
 END i177
 PIN i178
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 327.465 27.645 328.035 ;
  END
 END i178
 PIN i179
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 331.645 27.645 332.215 ;
  END
 END i179
 PIN i180
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 335.635 27.645 336.205 ;
  END
 END i180
 PIN i181
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 339.815 27.645 340.385 ;
  END
 END i181
 PIN i182
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 343.805 27.645 344.375 ;
  END
 END i182
 PIN i183
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 347.985 27.645 348.555 ;
  END
 END i183
 PIN i184
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 31.825 27.645 32.395 ;
  END
 END i184
 PIN i185
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 351.975 27.645 352.545 ;
  END
 END i185
 PIN i186
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 356.155 27.645 356.725 ;
  END
 END i186
 PIN i187
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 360.145 27.645 360.715 ;
  END
 END i187
 PIN i188
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 364.325 27.645 364.895 ;
  END
 END i188
 PIN i189
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 368.315 27.645 368.885 ;
  END
 END i189
 PIN i190
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 372.495 27.645 373.065 ;
  END
 END i190
 PIN i191
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 376.485 27.645 377.055 ;
  END
 END i191
 PIN i192
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 35.815 27.645 36.385 ;
  END
 END i192
 PIN i193
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 39.995 27.645 40.565 ;
  END
 END i193
 PIN i194
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 187.245 3.705 187.815 ;
  END
 END i194
 PIN i195
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 187.625 4.465 188.195 ;
  END
 END i195
 PIN i196
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 3.705 28.405 4.275 ;
  END
 END i196
 PIN i197
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 7.885 28.405 8.455 ;
  END
 END i197
 PIN i198
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 44.555 28.405 45.125 ;
  END
 END i198
 PIN i199
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 48.735 28.405 49.305 ;
  END
 END i199
 PIN i200
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 52.725 28.405 53.295 ;
  END
 END i200
 PIN i201
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 56.905 28.405 57.475 ;
  END
 END i201
 PIN i202
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 60.895 28.405 61.465 ;
  END
 END i202
 PIN i203
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 65.075 28.405 65.645 ;
  END
 END i203
 PIN i204
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 69.065 28.405 69.635 ;
  END
 END i204
 PIN i205
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 73.245 28.405 73.815 ;
  END
 END i205
 PIN i206
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 77.235 28.405 77.805 ;
  END
 END i206
 PIN i207
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 81.415 28.405 81.985 ;
  END
 END i207
 PIN i208
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 11.875 28.405 12.445 ;
  END
 END i208
 PIN i209
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 103.645 28.405 104.215 ;
  END
 END i209
 PIN i210
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 107.825 28.405 108.395 ;
  END
 END i210
 PIN i211
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 111.815 28.405 112.385 ;
  END
 END i211
 PIN i212
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 115.995 28.405 116.565 ;
  END
 END i212
 PIN i213
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 119.985 28.405 120.555 ;
  END
 END i213
 PIN i214
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 124.165 28.405 124.735 ;
  END
 END i214
 PIN i215
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 128.155 28.405 128.725 ;
  END
 END i215
 PIN i216
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 132.335 28.405 132.905 ;
  END
 END i216
 PIN i217
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 136.325 28.405 136.895 ;
  END
 END i217
 PIN i218
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 140.505 28.405 141.075 ;
  END
 END i218
 PIN i219
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 16.055 28.405 16.625 ;
  END
 END i219
 PIN i220
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 144.495 28.405 145.065 ;
  END
 END i220
 PIN i221
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 148.675 28.405 149.245 ;
  END
 END i221
 PIN i222
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 152.665 28.405 153.235 ;
  END
 END i222
 PIN i223
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 156.845 28.405 157.415 ;
  END
 END i223
 PIN i224
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 160.835 28.405 161.405 ;
  END
 END i224
 PIN i225
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 165.015 28.405 165.585 ;
  END
 END i225
 PIN i226
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 169.005 28.405 169.575 ;
  END
 END i226
 PIN i227
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 173.185 28.405 173.755 ;
  END
 END i227
 PIN i228
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 177.175 28.405 177.745 ;
  END
 END i228
 PIN i229
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 206.625 28.405 207.195 ;
  END
 END i229
 PIN i230
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 20.045 28.405 20.615 ;
  END
 END i230
 PIN i231
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 210.615 28.405 211.185 ;
  END
 END i231
 PIN i232
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 214.795 28.405 215.365 ;
  END
 END i232
 PIN i233
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 218.785 28.405 219.355 ;
  END
 END i233
 PIN i234
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 222.965 28.405 223.535 ;
  END
 END i234
 PIN i235
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 226.955 28.405 227.525 ;
  END
 END i235
 PIN i236
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 231.135 28.405 231.705 ;
  END
 END i236
 PIN i237
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 235.125 28.405 235.695 ;
  END
 END i237
 PIN i238
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 239.305 28.405 239.875 ;
  END
 END i238
 PIN i239
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 243.295 28.405 243.865 ;
  END
 END i239
 PIN i240
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 247.475 28.405 248.045 ;
  END
 END i240
 PIN i241
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 24.225 28.405 24.795 ;
  END
 END i241
 PIN i242
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 251.465 28.405 252.035 ;
  END
 END i242
 PIN i243
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 255.645 28.405 256.215 ;
  END
 END i243
 PIN i244
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 259.635 28.405 260.205 ;
  END
 END i244
 PIN i245
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 263.815 28.405 264.385 ;
  END
 END i245
 PIN i246
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 267.805 28.405 268.375 ;
  END
 END i246
 PIN i247
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 271.985 28.405 272.555 ;
  END
 END i247
 PIN i248
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 275.975 28.405 276.545 ;
  END
 END i248
 PIN i249
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 280.155 28.405 280.725 ;
  END
 END i249
 PIN i250
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 302.385 28.405 302.955 ;
  END
 END i250
 PIN i251
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 306.565 28.405 307.135 ;
  END
 END i251
 PIN i252
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 28.215 28.405 28.785 ;
  END
 END i252
 PIN i253
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 310.555 28.405 311.125 ;
  END
 END i253
 PIN i254
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 314.735 28.405 315.305 ;
  END
 END i254
 PIN i255
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 318.725 28.405 319.295 ;
  END
 END i255
 PIN i256
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 322.905 28.405 323.475 ;
  END
 END i256
 PIN i257
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 326.895 28.405 327.465 ;
  END
 END i257
 PIN i258
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 331.075 28.405 331.645 ;
  END
 END i258
 PIN i259
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 335.065 28.405 335.635 ;
  END
 END i259
 PIN i260
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 339.245 28.405 339.815 ;
  END
 END i260
 PIN i261
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 343.235 28.405 343.805 ;
  END
 END i261
 PIN i262
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 347.415 28.405 347.985 ;
  END
 END i262
 PIN i263
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 32.395 28.405 32.965 ;
  END
 END i263
 PIN i264
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 351.405 28.405 351.975 ;
  END
 END i264
 PIN i265
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 355.585 28.405 356.155 ;
  END
 END i265
 PIN i266
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 359.575 28.405 360.145 ;
  END
 END i266
 PIN i267
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 363.755 28.405 364.325 ;
  END
 END i267
 PIN i268
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 367.745 28.405 368.315 ;
  END
 END i268
 PIN i269
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 371.925 28.405 372.495 ;
  END
 END i269
 PIN i270
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 375.915 28.405 376.485 ;
  END
 END i270
 PIN i271
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 36.385 28.405 36.955 ;
  END
 END i271
 PIN i272
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 40.565 28.405 41.135 ;
  END
 END i272
 PIN i273
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 4.275 179.645 4.845 180.215 ;
  END
 END i273
 PIN i274
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 5.415 179.645 5.985 180.215 ;
  END
 END i274
 PIN i275
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 6.935 179.645 7.505 180.215 ;
  END
 END i275
 PIN i276
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 8.835 179.645 9.405 180.215 ;
  END
 END i276
 PIN i277
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 4.275 192.945 4.845 193.515 ;
  END
 END i277
 PIN i278
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 5.415 192.945 5.985 193.515 ;
  END
 END i278
 PIN i279
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 6.935 192.945 7.505 193.515 ;
  END
 END i279
 PIN i280
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 8.835 192.945 9.405 193.515 ;
  END
 END i280
 OBS
  LAYER metal1 ;
   RECT 23.18 0.0 157.32 1.71 ;
   RECT 23.18 1.71 157.32 3.42 ;
   RECT 23.18 3.42 157.32 5.13 ;
   RECT 23.18 5.13 157.32 6.84 ;
   RECT 23.18 6.84 157.32 8.55 ;
   RECT 23.18 8.55 157.32 10.26 ;
   RECT 23.18 10.26 157.32 11.97 ;
   RECT 23.18 11.97 157.32 13.68 ;
   RECT 23.18 13.68 157.32 15.39 ;
   RECT 23.18 15.39 157.32 17.1 ;
   RECT 23.18 17.1 157.32 18.81 ;
   RECT 23.18 18.81 157.32 20.52 ;
   RECT 23.18 20.52 157.32 22.23 ;
   RECT 23.18 22.23 157.32 23.94 ;
   RECT 23.18 23.94 157.32 25.65 ;
   RECT 23.18 25.65 157.32 27.36 ;
   RECT 23.18 27.36 157.32 29.07 ;
   RECT 23.18 29.07 157.32 30.78 ;
   RECT 23.18 30.78 157.32 32.49 ;
   RECT 23.18 32.49 157.32 34.2 ;
   RECT 23.18 34.2 157.32 35.91 ;
   RECT 23.18 35.91 157.32 37.62 ;
   RECT 23.18 37.62 157.32 39.33 ;
   RECT 23.18 39.33 157.32 41.04 ;
   RECT 23.18 41.04 157.32 42.75 ;
   RECT 23.18 42.75 157.32 44.46 ;
   RECT 23.18 44.46 157.32 46.17 ;
   RECT 23.18 46.17 157.32 47.88 ;
   RECT 23.18 47.88 157.32 49.59 ;
   RECT 23.18 49.59 157.32 51.3 ;
   RECT 23.18 51.3 157.32 53.01 ;
   RECT 23.18 53.01 157.32 54.72 ;
   RECT 23.18 54.72 157.32 56.43 ;
   RECT 23.18 56.43 157.32 58.14 ;
   RECT 23.18 58.14 157.32 59.85 ;
   RECT 23.18 59.85 157.32 61.56 ;
   RECT 23.18 61.56 157.32 63.27 ;
   RECT 23.18 63.27 157.32 64.98 ;
   RECT 23.18 64.98 157.32 66.69 ;
   RECT 23.18 66.69 157.32 68.4 ;
   RECT 23.18 68.4 157.32 70.11 ;
   RECT 23.18 70.11 157.32 71.82 ;
   RECT 23.18 71.82 157.32 73.53 ;
   RECT 23.18 73.53 157.32 75.24 ;
   RECT 23.18 75.24 157.32 76.95 ;
   RECT 23.18 76.95 157.32 78.66 ;
   RECT 23.18 78.66 157.32 80.37 ;
   RECT 23.18 80.37 157.32 82.08 ;
   RECT 23.18 82.08 157.32 83.79 ;
   RECT 23.18 83.79 157.32 85.5 ;
   RECT 23.18 85.5 157.32 87.21 ;
   RECT 23.18 87.21 157.32 88.92 ;
   RECT 23.18 88.92 157.32 90.63 ;
   RECT 23.18 90.63 157.32 92.34 ;
   RECT 23.18 92.34 157.32 94.05 ;
   RECT 23.18 94.05 157.32 95.76 ;
   RECT 23.18 95.76 157.32 97.47 ;
   RECT 23.18 97.47 157.32 99.18 ;
   RECT 23.18 99.18 157.32 100.89 ;
   RECT 23.18 100.89 157.32 102.6 ;
   RECT 23.18 102.6 157.32 104.31 ;
   RECT 23.18 104.31 157.32 106.02 ;
   RECT 23.18 106.02 157.32 107.73 ;
   RECT 23.18 107.73 157.32 109.44 ;
   RECT 23.18 109.44 157.32 111.15 ;
   RECT 23.18 111.15 157.32 112.86 ;
   RECT 23.18 112.86 157.32 114.57 ;
   RECT 23.18 114.57 157.32 116.28 ;
   RECT 23.18 116.28 157.32 117.99 ;
   RECT 23.18 117.99 157.32 119.7 ;
   RECT 23.18 119.7 157.32 121.41 ;
   RECT 23.18 121.41 157.32 123.12 ;
   RECT 23.18 123.12 157.32 124.83 ;
   RECT 23.18 124.83 157.32 126.54 ;
   RECT 23.18 126.54 157.32 128.25 ;
   RECT 23.18 128.25 157.32 129.96 ;
   RECT 23.18 129.96 157.32 131.67 ;
   RECT 23.18 131.67 157.32 133.38 ;
   RECT 23.18 133.38 157.32 135.09 ;
   RECT 23.18 135.09 157.32 136.8 ;
   RECT 23.18 136.8 157.32 138.51 ;
   RECT 23.18 138.51 157.32 140.22 ;
   RECT 23.18 140.22 157.32 141.93 ;
   RECT 23.18 141.93 157.32 143.64 ;
   RECT 23.18 143.64 157.32 145.35 ;
   RECT 23.18 145.35 157.32 147.06 ;
   RECT 23.18 147.06 157.32 148.77 ;
   RECT 23.18 148.77 157.32 150.48 ;
   RECT 23.18 150.48 157.32 152.19 ;
   RECT 23.18 152.19 157.32 153.9 ;
   RECT 23.18 153.9 157.32 155.61 ;
   RECT 23.18 155.61 157.32 157.32 ;
   RECT 23.18 157.32 157.32 159.03 ;
   RECT 23.18 159.03 157.32 160.74 ;
   RECT 23.18 160.74 157.32 162.45 ;
   RECT 23.18 162.45 157.32 164.16 ;
   RECT 23.18 164.16 157.32 165.87 ;
   RECT 23.18 165.87 157.32 167.58 ;
   RECT 23.18 167.58 157.32 169.29 ;
   RECT 23.18 169.29 157.32 171.0 ;
   RECT 23.18 171.0 157.32 172.71 ;
   RECT 23.18 172.71 157.32 174.42 ;
   RECT 23.18 174.42 157.32 176.13 ;
   RECT 23.18 176.13 157.32 177.84 ;
   RECT 0.0 177.84 157.32 179.55 ;
   RECT 0.0 179.55 157.32 181.26 ;
   RECT 0.0 181.26 157.32 182.97 ;
   RECT 0.0 182.97 157.32 184.68 ;
   RECT 0.0 184.68 157.32 186.39 ;
   RECT 0.0 186.39 157.32 188.1 ;
   RECT 0.0 188.1 157.32 189.81 ;
   RECT 0.0 189.81 157.32 191.52 ;
   RECT 0.0 191.52 157.32 193.23 ;
   RECT 0.0 193.23 157.32 194.94 ;
   RECT 0.0 194.94 157.32 196.65 ;
   RECT 0.0 196.65 157.32 198.36 ;
   RECT 0.0 198.36 157.32 200.07 ;
   RECT 0.0 200.07 157.32 201.78 ;
   RECT 0.0 201.78 157.32 203.49 ;
   RECT 0.0 203.49 157.32 205.2 ;
   RECT 0.0 205.2 157.32 206.91 ;
   RECT 23.18 206.91 157.32 208.62 ;
   RECT 23.18 208.62 157.32 210.33 ;
   RECT 23.18 210.33 157.32 212.04 ;
   RECT 23.18 212.04 157.32 213.75 ;
   RECT 23.18 213.75 157.32 215.46 ;
   RECT 23.18 215.46 157.32 217.17 ;
   RECT 23.18 217.17 157.32 218.88 ;
   RECT 23.18 218.88 157.32 220.59 ;
   RECT 23.18 220.59 157.32 222.3 ;
   RECT 23.18 222.3 157.32 224.01 ;
   RECT 23.18 224.01 157.32 225.72 ;
   RECT 23.18 225.72 157.32 227.43 ;
   RECT 23.18 227.43 157.32 229.14 ;
   RECT 23.18 229.14 157.32 230.85 ;
   RECT 23.18 230.85 157.32 232.56 ;
   RECT 23.18 232.56 157.32 234.27 ;
   RECT 23.18 234.27 157.32 235.98 ;
   RECT 23.18 235.98 157.32 237.69 ;
   RECT 23.18 237.69 157.32 239.4 ;
   RECT 23.18 239.4 157.32 241.11 ;
   RECT 23.18 241.11 157.32 242.82 ;
   RECT 23.18 242.82 157.32 244.53 ;
   RECT 23.18 244.53 157.32 246.24 ;
   RECT 23.18 246.24 157.32 247.95 ;
   RECT 23.18 247.95 157.32 249.66 ;
   RECT 23.18 249.66 157.32 251.37 ;
   RECT 23.18 251.37 157.32 253.08 ;
   RECT 23.18 253.08 157.32 254.79 ;
   RECT 23.18 254.79 157.32 256.5 ;
   RECT 23.18 256.5 157.32 258.21 ;
   RECT 23.18 258.21 157.32 259.92 ;
   RECT 23.18 259.92 157.32 261.63 ;
   RECT 23.18 261.63 157.32 263.34 ;
   RECT 23.18 263.34 157.32 265.05 ;
   RECT 23.18 265.05 157.32 266.76 ;
   RECT 23.18 266.76 157.32 268.47 ;
   RECT 23.18 268.47 157.32 270.18 ;
   RECT 23.18 270.18 157.32 271.89 ;
   RECT 23.18 271.89 157.32 273.6 ;
   RECT 23.18 273.6 157.32 275.31 ;
   RECT 23.18 275.31 157.32 277.02 ;
   RECT 23.18 277.02 157.32 278.73 ;
   RECT 23.18 278.73 157.32 280.44 ;
   RECT 23.18 280.44 157.32 282.15 ;
   RECT 23.18 282.15 157.32 283.86 ;
   RECT 23.18 283.86 157.32 285.57 ;
   RECT 23.18 285.57 157.32 287.28 ;
   RECT 23.18 287.28 157.32 288.99 ;
   RECT 23.18 288.99 157.32 290.7 ;
   RECT 23.18 290.7 157.32 292.41 ;
   RECT 23.18 292.41 157.32 294.12 ;
   RECT 23.18 294.12 157.32 295.83 ;
   RECT 23.18 295.83 157.32 297.54 ;
   RECT 23.18 297.54 157.32 299.25 ;
   RECT 23.18 299.25 157.32 300.96 ;
   RECT 23.18 300.96 157.32 302.67 ;
   RECT 23.18 302.67 157.32 304.38 ;
   RECT 23.18 304.38 157.32 306.09 ;
   RECT 23.18 306.09 157.32 307.8 ;
   RECT 23.18 307.8 157.32 309.51 ;
   RECT 23.18 309.51 157.32 311.22 ;
   RECT 23.18 311.22 157.32 312.93 ;
   RECT 23.18 312.93 157.32 314.64 ;
   RECT 23.18 314.64 157.32 316.35 ;
   RECT 23.18 316.35 157.32 318.06 ;
   RECT 23.18 318.06 157.32 319.77 ;
   RECT 23.18 319.77 157.32 321.48 ;
   RECT 23.18 321.48 157.32 323.19 ;
   RECT 23.18 323.19 157.32 324.9 ;
   RECT 23.18 324.9 157.32 326.61 ;
   RECT 23.18 326.61 157.32 328.32 ;
   RECT 23.18 328.32 157.32 330.03 ;
   RECT 23.18 330.03 157.32 331.74 ;
   RECT 23.18 331.74 157.32 333.45 ;
   RECT 23.18 333.45 157.32 335.16 ;
   RECT 23.18 335.16 157.32 336.87 ;
   RECT 23.18 336.87 157.32 338.58 ;
   RECT 23.18 338.58 157.32 340.29 ;
   RECT 23.18 340.29 157.32 342.0 ;
   RECT 23.18 342.0 157.32 343.71 ;
   RECT 23.18 343.71 157.32 345.42 ;
   RECT 23.18 345.42 157.32 347.13 ;
   RECT 23.18 347.13 157.32 348.84 ;
   RECT 23.18 348.84 157.32 350.55 ;
   RECT 23.18 350.55 157.32 352.26 ;
   RECT 23.18 352.26 157.32 353.97 ;
   RECT 23.18 353.97 157.32 355.68 ;
   RECT 23.18 355.68 157.32 357.39 ;
   RECT 23.18 357.39 157.32 359.1 ;
   RECT 23.18 359.1 157.32 360.81 ;
   RECT 23.18 360.81 157.32 362.52 ;
   RECT 23.18 362.52 157.32 364.23 ;
   RECT 23.18 364.23 157.32 365.94 ;
   RECT 23.18 365.94 157.32 367.65 ;
   RECT 23.18 367.65 157.32 369.36 ;
   RECT 23.18 369.36 157.32 371.07 ;
   RECT 23.18 371.07 157.32 372.78 ;
   RECT 23.18 372.78 157.32 374.49 ;
   RECT 23.18 374.49 157.32 376.2 ;
   RECT 23.18 376.2 157.32 377.91 ;
   RECT 23.18 377.91 157.32 379.62 ;
   RECT 23.18 379.62 157.32 381.33 ;
  LAYER via1 ;
   RECT 23.18 0.0 157.32 1.71 ;
   RECT 23.18 1.71 157.32 3.42 ;
   RECT 23.18 3.42 157.32 5.13 ;
   RECT 23.18 5.13 157.32 6.84 ;
   RECT 23.18 6.84 157.32 8.55 ;
   RECT 23.18 8.55 157.32 10.26 ;
   RECT 23.18 10.26 157.32 11.97 ;
   RECT 23.18 11.97 157.32 13.68 ;
   RECT 23.18 13.68 157.32 15.39 ;
   RECT 23.18 15.39 157.32 17.1 ;
   RECT 23.18 17.1 157.32 18.81 ;
   RECT 23.18 18.81 157.32 20.52 ;
   RECT 23.18 20.52 157.32 22.23 ;
   RECT 23.18 22.23 157.32 23.94 ;
   RECT 23.18 23.94 157.32 25.65 ;
   RECT 23.18 25.65 157.32 27.36 ;
   RECT 23.18 27.36 157.32 29.07 ;
   RECT 23.18 29.07 157.32 30.78 ;
   RECT 23.18 30.78 157.32 32.49 ;
   RECT 23.18 32.49 157.32 34.2 ;
   RECT 23.18 34.2 157.32 35.91 ;
   RECT 23.18 35.91 157.32 37.62 ;
   RECT 23.18 37.62 157.32 39.33 ;
   RECT 23.18 39.33 157.32 41.04 ;
   RECT 23.18 41.04 157.32 42.75 ;
   RECT 23.18 42.75 157.32 44.46 ;
   RECT 23.18 44.46 157.32 46.17 ;
   RECT 23.18 46.17 157.32 47.88 ;
   RECT 23.18 47.88 157.32 49.59 ;
   RECT 23.18 49.59 157.32 51.3 ;
   RECT 23.18 51.3 157.32 53.01 ;
   RECT 23.18 53.01 157.32 54.72 ;
   RECT 23.18 54.72 157.32 56.43 ;
   RECT 23.18 56.43 157.32 58.14 ;
   RECT 23.18 58.14 157.32 59.85 ;
   RECT 23.18 59.85 157.32 61.56 ;
   RECT 23.18 61.56 157.32 63.27 ;
   RECT 23.18 63.27 157.32 64.98 ;
   RECT 23.18 64.98 157.32 66.69 ;
   RECT 23.18 66.69 157.32 68.4 ;
   RECT 23.18 68.4 157.32 70.11 ;
   RECT 23.18 70.11 157.32 71.82 ;
   RECT 23.18 71.82 157.32 73.53 ;
   RECT 23.18 73.53 157.32 75.24 ;
   RECT 23.18 75.24 157.32 76.95 ;
   RECT 23.18 76.95 157.32 78.66 ;
   RECT 23.18 78.66 157.32 80.37 ;
   RECT 23.18 80.37 157.32 82.08 ;
   RECT 23.18 82.08 157.32 83.79 ;
   RECT 23.18 83.79 157.32 85.5 ;
   RECT 23.18 85.5 157.32 87.21 ;
   RECT 23.18 87.21 157.32 88.92 ;
   RECT 23.18 88.92 157.32 90.63 ;
   RECT 23.18 90.63 157.32 92.34 ;
   RECT 23.18 92.34 157.32 94.05 ;
   RECT 23.18 94.05 157.32 95.76 ;
   RECT 23.18 95.76 157.32 97.47 ;
   RECT 23.18 97.47 157.32 99.18 ;
   RECT 23.18 99.18 157.32 100.89 ;
   RECT 23.18 100.89 157.32 102.6 ;
   RECT 23.18 102.6 157.32 104.31 ;
   RECT 23.18 104.31 157.32 106.02 ;
   RECT 23.18 106.02 157.32 107.73 ;
   RECT 23.18 107.73 157.32 109.44 ;
   RECT 23.18 109.44 157.32 111.15 ;
   RECT 23.18 111.15 157.32 112.86 ;
   RECT 23.18 112.86 157.32 114.57 ;
   RECT 23.18 114.57 157.32 116.28 ;
   RECT 23.18 116.28 157.32 117.99 ;
   RECT 23.18 117.99 157.32 119.7 ;
   RECT 23.18 119.7 157.32 121.41 ;
   RECT 23.18 121.41 157.32 123.12 ;
   RECT 23.18 123.12 157.32 124.83 ;
   RECT 23.18 124.83 157.32 126.54 ;
   RECT 23.18 126.54 157.32 128.25 ;
   RECT 23.18 128.25 157.32 129.96 ;
   RECT 23.18 129.96 157.32 131.67 ;
   RECT 23.18 131.67 157.32 133.38 ;
   RECT 23.18 133.38 157.32 135.09 ;
   RECT 23.18 135.09 157.32 136.8 ;
   RECT 23.18 136.8 157.32 138.51 ;
   RECT 23.18 138.51 157.32 140.22 ;
   RECT 23.18 140.22 157.32 141.93 ;
   RECT 23.18 141.93 157.32 143.64 ;
   RECT 23.18 143.64 157.32 145.35 ;
   RECT 23.18 145.35 157.32 147.06 ;
   RECT 23.18 147.06 157.32 148.77 ;
   RECT 23.18 148.77 157.32 150.48 ;
   RECT 23.18 150.48 157.32 152.19 ;
   RECT 23.18 152.19 157.32 153.9 ;
   RECT 23.18 153.9 157.32 155.61 ;
   RECT 23.18 155.61 157.32 157.32 ;
   RECT 23.18 157.32 157.32 159.03 ;
   RECT 23.18 159.03 157.32 160.74 ;
   RECT 23.18 160.74 157.32 162.45 ;
   RECT 23.18 162.45 157.32 164.16 ;
   RECT 23.18 164.16 157.32 165.87 ;
   RECT 23.18 165.87 157.32 167.58 ;
   RECT 23.18 167.58 157.32 169.29 ;
   RECT 23.18 169.29 157.32 171.0 ;
   RECT 23.18 171.0 157.32 172.71 ;
   RECT 23.18 172.71 157.32 174.42 ;
   RECT 23.18 174.42 157.32 176.13 ;
   RECT 23.18 176.13 157.32 177.84 ;
   RECT 0.0 177.84 157.32 179.55 ;
   RECT 0.0 179.55 157.32 181.26 ;
   RECT 0.0 181.26 157.32 182.97 ;
   RECT 0.0 182.97 157.32 184.68 ;
   RECT 0.0 184.68 157.32 186.39 ;
   RECT 0.0 186.39 157.32 188.1 ;
   RECT 0.0 188.1 157.32 189.81 ;
   RECT 0.0 189.81 157.32 191.52 ;
   RECT 0.0 191.52 157.32 193.23 ;
   RECT 0.0 193.23 157.32 194.94 ;
   RECT 0.0 194.94 157.32 196.65 ;
   RECT 0.0 196.65 157.32 198.36 ;
   RECT 0.0 198.36 157.32 200.07 ;
   RECT 0.0 200.07 157.32 201.78 ;
   RECT 0.0 201.78 157.32 203.49 ;
   RECT 0.0 203.49 157.32 205.2 ;
   RECT 0.0 205.2 157.32 206.91 ;
   RECT 23.18 206.91 157.32 208.62 ;
   RECT 23.18 208.62 157.32 210.33 ;
   RECT 23.18 210.33 157.32 212.04 ;
   RECT 23.18 212.04 157.32 213.75 ;
   RECT 23.18 213.75 157.32 215.46 ;
   RECT 23.18 215.46 157.32 217.17 ;
   RECT 23.18 217.17 157.32 218.88 ;
   RECT 23.18 218.88 157.32 220.59 ;
   RECT 23.18 220.59 157.32 222.3 ;
   RECT 23.18 222.3 157.32 224.01 ;
   RECT 23.18 224.01 157.32 225.72 ;
   RECT 23.18 225.72 157.32 227.43 ;
   RECT 23.18 227.43 157.32 229.14 ;
   RECT 23.18 229.14 157.32 230.85 ;
   RECT 23.18 230.85 157.32 232.56 ;
   RECT 23.18 232.56 157.32 234.27 ;
   RECT 23.18 234.27 157.32 235.98 ;
   RECT 23.18 235.98 157.32 237.69 ;
   RECT 23.18 237.69 157.32 239.4 ;
   RECT 23.18 239.4 157.32 241.11 ;
   RECT 23.18 241.11 157.32 242.82 ;
   RECT 23.18 242.82 157.32 244.53 ;
   RECT 23.18 244.53 157.32 246.24 ;
   RECT 23.18 246.24 157.32 247.95 ;
   RECT 23.18 247.95 157.32 249.66 ;
   RECT 23.18 249.66 157.32 251.37 ;
   RECT 23.18 251.37 157.32 253.08 ;
   RECT 23.18 253.08 157.32 254.79 ;
   RECT 23.18 254.79 157.32 256.5 ;
   RECT 23.18 256.5 157.32 258.21 ;
   RECT 23.18 258.21 157.32 259.92 ;
   RECT 23.18 259.92 157.32 261.63 ;
   RECT 23.18 261.63 157.32 263.34 ;
   RECT 23.18 263.34 157.32 265.05 ;
   RECT 23.18 265.05 157.32 266.76 ;
   RECT 23.18 266.76 157.32 268.47 ;
   RECT 23.18 268.47 157.32 270.18 ;
   RECT 23.18 270.18 157.32 271.89 ;
   RECT 23.18 271.89 157.32 273.6 ;
   RECT 23.18 273.6 157.32 275.31 ;
   RECT 23.18 275.31 157.32 277.02 ;
   RECT 23.18 277.02 157.32 278.73 ;
   RECT 23.18 278.73 157.32 280.44 ;
   RECT 23.18 280.44 157.32 282.15 ;
   RECT 23.18 282.15 157.32 283.86 ;
   RECT 23.18 283.86 157.32 285.57 ;
   RECT 23.18 285.57 157.32 287.28 ;
   RECT 23.18 287.28 157.32 288.99 ;
   RECT 23.18 288.99 157.32 290.7 ;
   RECT 23.18 290.7 157.32 292.41 ;
   RECT 23.18 292.41 157.32 294.12 ;
   RECT 23.18 294.12 157.32 295.83 ;
   RECT 23.18 295.83 157.32 297.54 ;
   RECT 23.18 297.54 157.32 299.25 ;
   RECT 23.18 299.25 157.32 300.96 ;
   RECT 23.18 300.96 157.32 302.67 ;
   RECT 23.18 302.67 157.32 304.38 ;
   RECT 23.18 304.38 157.32 306.09 ;
   RECT 23.18 306.09 157.32 307.8 ;
   RECT 23.18 307.8 157.32 309.51 ;
   RECT 23.18 309.51 157.32 311.22 ;
   RECT 23.18 311.22 157.32 312.93 ;
   RECT 23.18 312.93 157.32 314.64 ;
   RECT 23.18 314.64 157.32 316.35 ;
   RECT 23.18 316.35 157.32 318.06 ;
   RECT 23.18 318.06 157.32 319.77 ;
   RECT 23.18 319.77 157.32 321.48 ;
   RECT 23.18 321.48 157.32 323.19 ;
   RECT 23.18 323.19 157.32 324.9 ;
   RECT 23.18 324.9 157.32 326.61 ;
   RECT 23.18 326.61 157.32 328.32 ;
   RECT 23.18 328.32 157.32 330.03 ;
   RECT 23.18 330.03 157.32 331.74 ;
   RECT 23.18 331.74 157.32 333.45 ;
   RECT 23.18 333.45 157.32 335.16 ;
   RECT 23.18 335.16 157.32 336.87 ;
   RECT 23.18 336.87 157.32 338.58 ;
   RECT 23.18 338.58 157.32 340.29 ;
   RECT 23.18 340.29 157.32 342.0 ;
   RECT 23.18 342.0 157.32 343.71 ;
   RECT 23.18 343.71 157.32 345.42 ;
   RECT 23.18 345.42 157.32 347.13 ;
   RECT 23.18 347.13 157.32 348.84 ;
   RECT 23.18 348.84 157.32 350.55 ;
   RECT 23.18 350.55 157.32 352.26 ;
   RECT 23.18 352.26 157.32 353.97 ;
   RECT 23.18 353.97 157.32 355.68 ;
   RECT 23.18 355.68 157.32 357.39 ;
   RECT 23.18 357.39 157.32 359.1 ;
   RECT 23.18 359.1 157.32 360.81 ;
   RECT 23.18 360.81 157.32 362.52 ;
   RECT 23.18 362.52 157.32 364.23 ;
   RECT 23.18 364.23 157.32 365.94 ;
   RECT 23.18 365.94 157.32 367.65 ;
   RECT 23.18 367.65 157.32 369.36 ;
   RECT 23.18 369.36 157.32 371.07 ;
   RECT 23.18 371.07 157.32 372.78 ;
   RECT 23.18 372.78 157.32 374.49 ;
   RECT 23.18 374.49 157.32 376.2 ;
   RECT 23.18 376.2 157.32 377.91 ;
   RECT 23.18 377.91 157.32 379.62 ;
   RECT 23.18 379.62 157.32 381.33 ;
  LAYER metal2 ;
   RECT 23.18 0.0 157.32 1.71 ;
   RECT 23.18 1.71 157.32 3.42 ;
   RECT 23.18 3.42 157.32 5.13 ;
   RECT 23.18 5.13 157.32 6.84 ;
   RECT 23.18 6.84 157.32 8.55 ;
   RECT 23.18 8.55 157.32 10.26 ;
   RECT 23.18 10.26 157.32 11.97 ;
   RECT 23.18 11.97 157.32 13.68 ;
   RECT 23.18 13.68 157.32 15.39 ;
   RECT 23.18 15.39 157.32 17.1 ;
   RECT 23.18 17.1 157.32 18.81 ;
   RECT 23.18 18.81 157.32 20.52 ;
   RECT 23.18 20.52 157.32 22.23 ;
   RECT 23.18 22.23 157.32 23.94 ;
   RECT 23.18 23.94 157.32 25.65 ;
   RECT 23.18 25.65 157.32 27.36 ;
   RECT 23.18 27.36 157.32 29.07 ;
   RECT 23.18 29.07 157.32 30.78 ;
   RECT 23.18 30.78 157.32 32.49 ;
   RECT 23.18 32.49 157.32 34.2 ;
   RECT 23.18 34.2 157.32 35.91 ;
   RECT 23.18 35.91 157.32 37.62 ;
   RECT 23.18 37.62 157.32 39.33 ;
   RECT 23.18 39.33 157.32 41.04 ;
   RECT 23.18 41.04 157.32 42.75 ;
   RECT 23.18 42.75 157.32 44.46 ;
   RECT 23.18 44.46 157.32 46.17 ;
   RECT 23.18 46.17 157.32 47.88 ;
   RECT 23.18 47.88 157.32 49.59 ;
   RECT 23.18 49.59 157.32 51.3 ;
   RECT 23.18 51.3 157.32 53.01 ;
   RECT 23.18 53.01 157.32 54.72 ;
   RECT 23.18 54.72 157.32 56.43 ;
   RECT 23.18 56.43 157.32 58.14 ;
   RECT 23.18 58.14 157.32 59.85 ;
   RECT 23.18 59.85 157.32 61.56 ;
   RECT 23.18 61.56 157.32 63.27 ;
   RECT 23.18 63.27 157.32 64.98 ;
   RECT 23.18 64.98 157.32 66.69 ;
   RECT 23.18 66.69 157.32 68.4 ;
   RECT 23.18 68.4 157.32 70.11 ;
   RECT 23.18 70.11 157.32 71.82 ;
   RECT 23.18 71.82 157.32 73.53 ;
   RECT 23.18 73.53 157.32 75.24 ;
   RECT 23.18 75.24 157.32 76.95 ;
   RECT 23.18 76.95 157.32 78.66 ;
   RECT 23.18 78.66 157.32 80.37 ;
   RECT 23.18 80.37 157.32 82.08 ;
   RECT 23.18 82.08 157.32 83.79 ;
   RECT 23.18 83.79 157.32 85.5 ;
   RECT 23.18 85.5 157.32 87.21 ;
   RECT 23.18 87.21 157.32 88.92 ;
   RECT 23.18 88.92 157.32 90.63 ;
   RECT 23.18 90.63 157.32 92.34 ;
   RECT 23.18 92.34 157.32 94.05 ;
   RECT 23.18 94.05 157.32 95.76 ;
   RECT 23.18 95.76 157.32 97.47 ;
   RECT 23.18 97.47 157.32 99.18 ;
   RECT 23.18 99.18 157.32 100.89 ;
   RECT 23.18 100.89 157.32 102.6 ;
   RECT 23.18 102.6 157.32 104.31 ;
   RECT 23.18 104.31 157.32 106.02 ;
   RECT 23.18 106.02 157.32 107.73 ;
   RECT 23.18 107.73 157.32 109.44 ;
   RECT 23.18 109.44 157.32 111.15 ;
   RECT 23.18 111.15 157.32 112.86 ;
   RECT 23.18 112.86 157.32 114.57 ;
   RECT 23.18 114.57 157.32 116.28 ;
   RECT 23.18 116.28 157.32 117.99 ;
   RECT 23.18 117.99 157.32 119.7 ;
   RECT 23.18 119.7 157.32 121.41 ;
   RECT 23.18 121.41 157.32 123.12 ;
   RECT 23.18 123.12 157.32 124.83 ;
   RECT 23.18 124.83 157.32 126.54 ;
   RECT 23.18 126.54 157.32 128.25 ;
   RECT 23.18 128.25 157.32 129.96 ;
   RECT 23.18 129.96 157.32 131.67 ;
   RECT 23.18 131.67 157.32 133.38 ;
   RECT 23.18 133.38 157.32 135.09 ;
   RECT 23.18 135.09 157.32 136.8 ;
   RECT 23.18 136.8 157.32 138.51 ;
   RECT 23.18 138.51 157.32 140.22 ;
   RECT 23.18 140.22 157.32 141.93 ;
   RECT 23.18 141.93 157.32 143.64 ;
   RECT 23.18 143.64 157.32 145.35 ;
   RECT 23.18 145.35 157.32 147.06 ;
   RECT 23.18 147.06 157.32 148.77 ;
   RECT 23.18 148.77 157.32 150.48 ;
   RECT 23.18 150.48 157.32 152.19 ;
   RECT 23.18 152.19 157.32 153.9 ;
   RECT 23.18 153.9 157.32 155.61 ;
   RECT 23.18 155.61 157.32 157.32 ;
   RECT 23.18 157.32 157.32 159.03 ;
   RECT 23.18 159.03 157.32 160.74 ;
   RECT 23.18 160.74 157.32 162.45 ;
   RECT 23.18 162.45 157.32 164.16 ;
   RECT 23.18 164.16 157.32 165.87 ;
   RECT 23.18 165.87 157.32 167.58 ;
   RECT 23.18 167.58 157.32 169.29 ;
   RECT 23.18 169.29 157.32 171.0 ;
   RECT 23.18 171.0 157.32 172.71 ;
   RECT 23.18 172.71 157.32 174.42 ;
   RECT 23.18 174.42 157.32 176.13 ;
   RECT 23.18 176.13 157.32 177.84 ;
   RECT 0.0 177.84 157.32 179.55 ;
   RECT 0.0 179.55 157.32 181.26 ;
   RECT 0.0 181.26 157.32 182.97 ;
   RECT 0.0 182.97 157.32 184.68 ;
   RECT 0.0 184.68 157.32 186.39 ;
   RECT 0.0 186.39 157.32 188.1 ;
   RECT 0.0 188.1 157.32 189.81 ;
   RECT 0.0 189.81 157.32 191.52 ;
   RECT 0.0 191.52 157.32 193.23 ;
   RECT 0.0 193.23 157.32 194.94 ;
   RECT 0.0 194.94 157.32 196.65 ;
   RECT 0.0 196.65 157.32 198.36 ;
   RECT 0.0 198.36 157.32 200.07 ;
   RECT 0.0 200.07 157.32 201.78 ;
   RECT 0.0 201.78 157.32 203.49 ;
   RECT 0.0 203.49 157.32 205.2 ;
   RECT 0.0 205.2 157.32 206.91 ;
   RECT 23.18 206.91 157.32 208.62 ;
   RECT 23.18 208.62 157.32 210.33 ;
   RECT 23.18 210.33 157.32 212.04 ;
   RECT 23.18 212.04 157.32 213.75 ;
   RECT 23.18 213.75 157.32 215.46 ;
   RECT 23.18 215.46 157.32 217.17 ;
   RECT 23.18 217.17 157.32 218.88 ;
   RECT 23.18 218.88 157.32 220.59 ;
   RECT 23.18 220.59 157.32 222.3 ;
   RECT 23.18 222.3 157.32 224.01 ;
   RECT 23.18 224.01 157.32 225.72 ;
   RECT 23.18 225.72 157.32 227.43 ;
   RECT 23.18 227.43 157.32 229.14 ;
   RECT 23.18 229.14 157.32 230.85 ;
   RECT 23.18 230.85 157.32 232.56 ;
   RECT 23.18 232.56 157.32 234.27 ;
   RECT 23.18 234.27 157.32 235.98 ;
   RECT 23.18 235.98 157.32 237.69 ;
   RECT 23.18 237.69 157.32 239.4 ;
   RECT 23.18 239.4 157.32 241.11 ;
   RECT 23.18 241.11 157.32 242.82 ;
   RECT 23.18 242.82 157.32 244.53 ;
   RECT 23.18 244.53 157.32 246.24 ;
   RECT 23.18 246.24 157.32 247.95 ;
   RECT 23.18 247.95 157.32 249.66 ;
   RECT 23.18 249.66 157.32 251.37 ;
   RECT 23.18 251.37 157.32 253.08 ;
   RECT 23.18 253.08 157.32 254.79 ;
   RECT 23.18 254.79 157.32 256.5 ;
   RECT 23.18 256.5 157.32 258.21 ;
   RECT 23.18 258.21 157.32 259.92 ;
   RECT 23.18 259.92 157.32 261.63 ;
   RECT 23.18 261.63 157.32 263.34 ;
   RECT 23.18 263.34 157.32 265.05 ;
   RECT 23.18 265.05 157.32 266.76 ;
   RECT 23.18 266.76 157.32 268.47 ;
   RECT 23.18 268.47 157.32 270.18 ;
   RECT 23.18 270.18 157.32 271.89 ;
   RECT 23.18 271.89 157.32 273.6 ;
   RECT 23.18 273.6 157.32 275.31 ;
   RECT 23.18 275.31 157.32 277.02 ;
   RECT 23.18 277.02 157.32 278.73 ;
   RECT 23.18 278.73 157.32 280.44 ;
   RECT 23.18 280.44 157.32 282.15 ;
   RECT 23.18 282.15 157.32 283.86 ;
   RECT 23.18 283.86 157.32 285.57 ;
   RECT 23.18 285.57 157.32 287.28 ;
   RECT 23.18 287.28 157.32 288.99 ;
   RECT 23.18 288.99 157.32 290.7 ;
   RECT 23.18 290.7 157.32 292.41 ;
   RECT 23.18 292.41 157.32 294.12 ;
   RECT 23.18 294.12 157.32 295.83 ;
   RECT 23.18 295.83 157.32 297.54 ;
   RECT 23.18 297.54 157.32 299.25 ;
   RECT 23.18 299.25 157.32 300.96 ;
   RECT 23.18 300.96 157.32 302.67 ;
   RECT 23.18 302.67 157.32 304.38 ;
   RECT 23.18 304.38 157.32 306.09 ;
   RECT 23.18 306.09 157.32 307.8 ;
   RECT 23.18 307.8 157.32 309.51 ;
   RECT 23.18 309.51 157.32 311.22 ;
   RECT 23.18 311.22 157.32 312.93 ;
   RECT 23.18 312.93 157.32 314.64 ;
   RECT 23.18 314.64 157.32 316.35 ;
   RECT 23.18 316.35 157.32 318.06 ;
   RECT 23.18 318.06 157.32 319.77 ;
   RECT 23.18 319.77 157.32 321.48 ;
   RECT 23.18 321.48 157.32 323.19 ;
   RECT 23.18 323.19 157.32 324.9 ;
   RECT 23.18 324.9 157.32 326.61 ;
   RECT 23.18 326.61 157.32 328.32 ;
   RECT 23.18 328.32 157.32 330.03 ;
   RECT 23.18 330.03 157.32 331.74 ;
   RECT 23.18 331.74 157.32 333.45 ;
   RECT 23.18 333.45 157.32 335.16 ;
   RECT 23.18 335.16 157.32 336.87 ;
   RECT 23.18 336.87 157.32 338.58 ;
   RECT 23.18 338.58 157.32 340.29 ;
   RECT 23.18 340.29 157.32 342.0 ;
   RECT 23.18 342.0 157.32 343.71 ;
   RECT 23.18 343.71 157.32 345.42 ;
   RECT 23.18 345.42 157.32 347.13 ;
   RECT 23.18 347.13 157.32 348.84 ;
   RECT 23.18 348.84 157.32 350.55 ;
   RECT 23.18 350.55 157.32 352.26 ;
   RECT 23.18 352.26 157.32 353.97 ;
   RECT 23.18 353.97 157.32 355.68 ;
   RECT 23.18 355.68 157.32 357.39 ;
   RECT 23.18 357.39 157.32 359.1 ;
   RECT 23.18 359.1 157.32 360.81 ;
   RECT 23.18 360.81 157.32 362.52 ;
   RECT 23.18 362.52 157.32 364.23 ;
   RECT 23.18 364.23 157.32 365.94 ;
   RECT 23.18 365.94 157.32 367.65 ;
   RECT 23.18 367.65 157.32 369.36 ;
   RECT 23.18 369.36 157.32 371.07 ;
   RECT 23.18 371.07 157.32 372.78 ;
   RECT 23.18 372.78 157.32 374.49 ;
   RECT 23.18 374.49 157.32 376.2 ;
   RECT 23.18 376.2 157.32 377.91 ;
   RECT 23.18 377.91 157.32 379.62 ;
   RECT 23.18 379.62 157.32 381.33 ;
  LAYER via2 ;
   RECT 23.18 0.0 157.32 1.71 ;
   RECT 23.18 1.71 157.32 3.42 ;
   RECT 23.18 3.42 157.32 5.13 ;
   RECT 23.18 5.13 157.32 6.84 ;
   RECT 23.18 6.84 157.32 8.55 ;
   RECT 23.18 8.55 157.32 10.26 ;
   RECT 23.18 10.26 157.32 11.97 ;
   RECT 23.18 11.97 157.32 13.68 ;
   RECT 23.18 13.68 157.32 15.39 ;
   RECT 23.18 15.39 157.32 17.1 ;
   RECT 23.18 17.1 157.32 18.81 ;
   RECT 23.18 18.81 157.32 20.52 ;
   RECT 23.18 20.52 157.32 22.23 ;
   RECT 23.18 22.23 157.32 23.94 ;
   RECT 23.18 23.94 157.32 25.65 ;
   RECT 23.18 25.65 157.32 27.36 ;
   RECT 23.18 27.36 157.32 29.07 ;
   RECT 23.18 29.07 157.32 30.78 ;
   RECT 23.18 30.78 157.32 32.49 ;
   RECT 23.18 32.49 157.32 34.2 ;
   RECT 23.18 34.2 157.32 35.91 ;
   RECT 23.18 35.91 157.32 37.62 ;
   RECT 23.18 37.62 157.32 39.33 ;
   RECT 23.18 39.33 157.32 41.04 ;
   RECT 23.18 41.04 157.32 42.75 ;
   RECT 23.18 42.75 157.32 44.46 ;
   RECT 23.18 44.46 157.32 46.17 ;
   RECT 23.18 46.17 157.32 47.88 ;
   RECT 23.18 47.88 157.32 49.59 ;
   RECT 23.18 49.59 157.32 51.3 ;
   RECT 23.18 51.3 157.32 53.01 ;
   RECT 23.18 53.01 157.32 54.72 ;
   RECT 23.18 54.72 157.32 56.43 ;
   RECT 23.18 56.43 157.32 58.14 ;
   RECT 23.18 58.14 157.32 59.85 ;
   RECT 23.18 59.85 157.32 61.56 ;
   RECT 23.18 61.56 157.32 63.27 ;
   RECT 23.18 63.27 157.32 64.98 ;
   RECT 23.18 64.98 157.32 66.69 ;
   RECT 23.18 66.69 157.32 68.4 ;
   RECT 23.18 68.4 157.32 70.11 ;
   RECT 23.18 70.11 157.32 71.82 ;
   RECT 23.18 71.82 157.32 73.53 ;
   RECT 23.18 73.53 157.32 75.24 ;
   RECT 23.18 75.24 157.32 76.95 ;
   RECT 23.18 76.95 157.32 78.66 ;
   RECT 23.18 78.66 157.32 80.37 ;
   RECT 23.18 80.37 157.32 82.08 ;
   RECT 23.18 82.08 157.32 83.79 ;
   RECT 23.18 83.79 157.32 85.5 ;
   RECT 23.18 85.5 157.32 87.21 ;
   RECT 23.18 87.21 157.32 88.92 ;
   RECT 23.18 88.92 157.32 90.63 ;
   RECT 23.18 90.63 157.32 92.34 ;
   RECT 23.18 92.34 157.32 94.05 ;
   RECT 23.18 94.05 157.32 95.76 ;
   RECT 23.18 95.76 157.32 97.47 ;
   RECT 23.18 97.47 157.32 99.18 ;
   RECT 23.18 99.18 157.32 100.89 ;
   RECT 23.18 100.89 157.32 102.6 ;
   RECT 23.18 102.6 157.32 104.31 ;
   RECT 23.18 104.31 157.32 106.02 ;
   RECT 23.18 106.02 157.32 107.73 ;
   RECT 23.18 107.73 157.32 109.44 ;
   RECT 23.18 109.44 157.32 111.15 ;
   RECT 23.18 111.15 157.32 112.86 ;
   RECT 23.18 112.86 157.32 114.57 ;
   RECT 23.18 114.57 157.32 116.28 ;
   RECT 23.18 116.28 157.32 117.99 ;
   RECT 23.18 117.99 157.32 119.7 ;
   RECT 23.18 119.7 157.32 121.41 ;
   RECT 23.18 121.41 157.32 123.12 ;
   RECT 23.18 123.12 157.32 124.83 ;
   RECT 23.18 124.83 157.32 126.54 ;
   RECT 23.18 126.54 157.32 128.25 ;
   RECT 23.18 128.25 157.32 129.96 ;
   RECT 23.18 129.96 157.32 131.67 ;
   RECT 23.18 131.67 157.32 133.38 ;
   RECT 23.18 133.38 157.32 135.09 ;
   RECT 23.18 135.09 157.32 136.8 ;
   RECT 23.18 136.8 157.32 138.51 ;
   RECT 23.18 138.51 157.32 140.22 ;
   RECT 23.18 140.22 157.32 141.93 ;
   RECT 23.18 141.93 157.32 143.64 ;
   RECT 23.18 143.64 157.32 145.35 ;
   RECT 23.18 145.35 157.32 147.06 ;
   RECT 23.18 147.06 157.32 148.77 ;
   RECT 23.18 148.77 157.32 150.48 ;
   RECT 23.18 150.48 157.32 152.19 ;
   RECT 23.18 152.19 157.32 153.9 ;
   RECT 23.18 153.9 157.32 155.61 ;
   RECT 23.18 155.61 157.32 157.32 ;
   RECT 23.18 157.32 157.32 159.03 ;
   RECT 23.18 159.03 157.32 160.74 ;
   RECT 23.18 160.74 157.32 162.45 ;
   RECT 23.18 162.45 157.32 164.16 ;
   RECT 23.18 164.16 157.32 165.87 ;
   RECT 23.18 165.87 157.32 167.58 ;
   RECT 23.18 167.58 157.32 169.29 ;
   RECT 23.18 169.29 157.32 171.0 ;
   RECT 23.18 171.0 157.32 172.71 ;
   RECT 23.18 172.71 157.32 174.42 ;
   RECT 23.18 174.42 157.32 176.13 ;
   RECT 23.18 176.13 157.32 177.84 ;
   RECT 0.0 177.84 157.32 179.55 ;
   RECT 0.0 179.55 157.32 181.26 ;
   RECT 0.0 181.26 157.32 182.97 ;
   RECT 0.0 182.97 157.32 184.68 ;
   RECT 0.0 184.68 157.32 186.39 ;
   RECT 0.0 186.39 157.32 188.1 ;
   RECT 0.0 188.1 157.32 189.81 ;
   RECT 0.0 189.81 157.32 191.52 ;
   RECT 0.0 191.52 157.32 193.23 ;
   RECT 0.0 193.23 157.32 194.94 ;
   RECT 0.0 194.94 157.32 196.65 ;
   RECT 0.0 196.65 157.32 198.36 ;
   RECT 0.0 198.36 157.32 200.07 ;
   RECT 0.0 200.07 157.32 201.78 ;
   RECT 0.0 201.78 157.32 203.49 ;
   RECT 0.0 203.49 157.32 205.2 ;
   RECT 0.0 205.2 157.32 206.91 ;
   RECT 23.18 206.91 157.32 208.62 ;
   RECT 23.18 208.62 157.32 210.33 ;
   RECT 23.18 210.33 157.32 212.04 ;
   RECT 23.18 212.04 157.32 213.75 ;
   RECT 23.18 213.75 157.32 215.46 ;
   RECT 23.18 215.46 157.32 217.17 ;
   RECT 23.18 217.17 157.32 218.88 ;
   RECT 23.18 218.88 157.32 220.59 ;
   RECT 23.18 220.59 157.32 222.3 ;
   RECT 23.18 222.3 157.32 224.01 ;
   RECT 23.18 224.01 157.32 225.72 ;
   RECT 23.18 225.72 157.32 227.43 ;
   RECT 23.18 227.43 157.32 229.14 ;
   RECT 23.18 229.14 157.32 230.85 ;
   RECT 23.18 230.85 157.32 232.56 ;
   RECT 23.18 232.56 157.32 234.27 ;
   RECT 23.18 234.27 157.32 235.98 ;
   RECT 23.18 235.98 157.32 237.69 ;
   RECT 23.18 237.69 157.32 239.4 ;
   RECT 23.18 239.4 157.32 241.11 ;
   RECT 23.18 241.11 157.32 242.82 ;
   RECT 23.18 242.82 157.32 244.53 ;
   RECT 23.18 244.53 157.32 246.24 ;
   RECT 23.18 246.24 157.32 247.95 ;
   RECT 23.18 247.95 157.32 249.66 ;
   RECT 23.18 249.66 157.32 251.37 ;
   RECT 23.18 251.37 157.32 253.08 ;
   RECT 23.18 253.08 157.32 254.79 ;
   RECT 23.18 254.79 157.32 256.5 ;
   RECT 23.18 256.5 157.32 258.21 ;
   RECT 23.18 258.21 157.32 259.92 ;
   RECT 23.18 259.92 157.32 261.63 ;
   RECT 23.18 261.63 157.32 263.34 ;
   RECT 23.18 263.34 157.32 265.05 ;
   RECT 23.18 265.05 157.32 266.76 ;
   RECT 23.18 266.76 157.32 268.47 ;
   RECT 23.18 268.47 157.32 270.18 ;
   RECT 23.18 270.18 157.32 271.89 ;
   RECT 23.18 271.89 157.32 273.6 ;
   RECT 23.18 273.6 157.32 275.31 ;
   RECT 23.18 275.31 157.32 277.02 ;
   RECT 23.18 277.02 157.32 278.73 ;
   RECT 23.18 278.73 157.32 280.44 ;
   RECT 23.18 280.44 157.32 282.15 ;
   RECT 23.18 282.15 157.32 283.86 ;
   RECT 23.18 283.86 157.32 285.57 ;
   RECT 23.18 285.57 157.32 287.28 ;
   RECT 23.18 287.28 157.32 288.99 ;
   RECT 23.18 288.99 157.32 290.7 ;
   RECT 23.18 290.7 157.32 292.41 ;
   RECT 23.18 292.41 157.32 294.12 ;
   RECT 23.18 294.12 157.32 295.83 ;
   RECT 23.18 295.83 157.32 297.54 ;
   RECT 23.18 297.54 157.32 299.25 ;
   RECT 23.18 299.25 157.32 300.96 ;
   RECT 23.18 300.96 157.32 302.67 ;
   RECT 23.18 302.67 157.32 304.38 ;
   RECT 23.18 304.38 157.32 306.09 ;
   RECT 23.18 306.09 157.32 307.8 ;
   RECT 23.18 307.8 157.32 309.51 ;
   RECT 23.18 309.51 157.32 311.22 ;
   RECT 23.18 311.22 157.32 312.93 ;
   RECT 23.18 312.93 157.32 314.64 ;
   RECT 23.18 314.64 157.32 316.35 ;
   RECT 23.18 316.35 157.32 318.06 ;
   RECT 23.18 318.06 157.32 319.77 ;
   RECT 23.18 319.77 157.32 321.48 ;
   RECT 23.18 321.48 157.32 323.19 ;
   RECT 23.18 323.19 157.32 324.9 ;
   RECT 23.18 324.9 157.32 326.61 ;
   RECT 23.18 326.61 157.32 328.32 ;
   RECT 23.18 328.32 157.32 330.03 ;
   RECT 23.18 330.03 157.32 331.74 ;
   RECT 23.18 331.74 157.32 333.45 ;
   RECT 23.18 333.45 157.32 335.16 ;
   RECT 23.18 335.16 157.32 336.87 ;
   RECT 23.18 336.87 157.32 338.58 ;
   RECT 23.18 338.58 157.32 340.29 ;
   RECT 23.18 340.29 157.32 342.0 ;
   RECT 23.18 342.0 157.32 343.71 ;
   RECT 23.18 343.71 157.32 345.42 ;
   RECT 23.18 345.42 157.32 347.13 ;
   RECT 23.18 347.13 157.32 348.84 ;
   RECT 23.18 348.84 157.32 350.55 ;
   RECT 23.18 350.55 157.32 352.26 ;
   RECT 23.18 352.26 157.32 353.97 ;
   RECT 23.18 353.97 157.32 355.68 ;
   RECT 23.18 355.68 157.32 357.39 ;
   RECT 23.18 357.39 157.32 359.1 ;
   RECT 23.18 359.1 157.32 360.81 ;
   RECT 23.18 360.81 157.32 362.52 ;
   RECT 23.18 362.52 157.32 364.23 ;
   RECT 23.18 364.23 157.32 365.94 ;
   RECT 23.18 365.94 157.32 367.65 ;
   RECT 23.18 367.65 157.32 369.36 ;
   RECT 23.18 369.36 157.32 371.07 ;
   RECT 23.18 371.07 157.32 372.78 ;
   RECT 23.18 372.78 157.32 374.49 ;
   RECT 23.18 374.49 157.32 376.2 ;
   RECT 23.18 376.2 157.32 377.91 ;
   RECT 23.18 377.91 157.32 379.62 ;
   RECT 23.18 379.62 157.32 381.33 ;
  LAYER metal3 ;
   RECT 23.18 0.0 157.32 1.71 ;
   RECT 23.18 1.71 157.32 3.42 ;
   RECT 23.18 3.42 157.32 5.13 ;
   RECT 23.18 5.13 157.32 6.84 ;
   RECT 23.18 6.84 157.32 8.55 ;
   RECT 23.18 8.55 157.32 10.26 ;
   RECT 23.18 10.26 157.32 11.97 ;
   RECT 23.18 11.97 157.32 13.68 ;
   RECT 23.18 13.68 157.32 15.39 ;
   RECT 23.18 15.39 157.32 17.1 ;
   RECT 23.18 17.1 157.32 18.81 ;
   RECT 23.18 18.81 157.32 20.52 ;
   RECT 23.18 20.52 157.32 22.23 ;
   RECT 23.18 22.23 157.32 23.94 ;
   RECT 23.18 23.94 157.32 25.65 ;
   RECT 23.18 25.65 157.32 27.36 ;
   RECT 23.18 27.36 157.32 29.07 ;
   RECT 23.18 29.07 157.32 30.78 ;
   RECT 23.18 30.78 157.32 32.49 ;
   RECT 23.18 32.49 157.32 34.2 ;
   RECT 23.18 34.2 157.32 35.91 ;
   RECT 23.18 35.91 157.32 37.62 ;
   RECT 23.18 37.62 157.32 39.33 ;
   RECT 23.18 39.33 157.32 41.04 ;
   RECT 23.18 41.04 157.32 42.75 ;
   RECT 23.18 42.75 157.32 44.46 ;
   RECT 23.18 44.46 157.32 46.17 ;
   RECT 23.18 46.17 157.32 47.88 ;
   RECT 23.18 47.88 157.32 49.59 ;
   RECT 23.18 49.59 157.32 51.3 ;
   RECT 23.18 51.3 157.32 53.01 ;
   RECT 23.18 53.01 157.32 54.72 ;
   RECT 23.18 54.72 157.32 56.43 ;
   RECT 23.18 56.43 157.32 58.14 ;
   RECT 23.18 58.14 157.32 59.85 ;
   RECT 23.18 59.85 157.32 61.56 ;
   RECT 23.18 61.56 157.32 63.27 ;
   RECT 23.18 63.27 157.32 64.98 ;
   RECT 23.18 64.98 157.32 66.69 ;
   RECT 23.18 66.69 157.32 68.4 ;
   RECT 23.18 68.4 157.32 70.11 ;
   RECT 23.18 70.11 157.32 71.82 ;
   RECT 23.18 71.82 157.32 73.53 ;
   RECT 23.18 73.53 157.32 75.24 ;
   RECT 23.18 75.24 157.32 76.95 ;
   RECT 23.18 76.95 157.32 78.66 ;
   RECT 23.18 78.66 157.32 80.37 ;
   RECT 23.18 80.37 157.32 82.08 ;
   RECT 23.18 82.08 157.32 83.79 ;
   RECT 23.18 83.79 157.32 85.5 ;
   RECT 23.18 85.5 157.32 87.21 ;
   RECT 23.18 87.21 157.32 88.92 ;
   RECT 23.18 88.92 157.32 90.63 ;
   RECT 23.18 90.63 157.32 92.34 ;
   RECT 23.18 92.34 157.32 94.05 ;
   RECT 23.18 94.05 157.32 95.76 ;
   RECT 23.18 95.76 157.32 97.47 ;
   RECT 23.18 97.47 157.32 99.18 ;
   RECT 23.18 99.18 157.32 100.89 ;
   RECT 23.18 100.89 157.32 102.6 ;
   RECT 23.18 102.6 157.32 104.31 ;
   RECT 23.18 104.31 157.32 106.02 ;
   RECT 23.18 106.02 157.32 107.73 ;
   RECT 23.18 107.73 157.32 109.44 ;
   RECT 23.18 109.44 157.32 111.15 ;
   RECT 23.18 111.15 157.32 112.86 ;
   RECT 23.18 112.86 157.32 114.57 ;
   RECT 23.18 114.57 157.32 116.28 ;
   RECT 23.18 116.28 157.32 117.99 ;
   RECT 23.18 117.99 157.32 119.7 ;
   RECT 23.18 119.7 157.32 121.41 ;
   RECT 23.18 121.41 157.32 123.12 ;
   RECT 23.18 123.12 157.32 124.83 ;
   RECT 23.18 124.83 157.32 126.54 ;
   RECT 23.18 126.54 157.32 128.25 ;
   RECT 23.18 128.25 157.32 129.96 ;
   RECT 23.18 129.96 157.32 131.67 ;
   RECT 23.18 131.67 157.32 133.38 ;
   RECT 23.18 133.38 157.32 135.09 ;
   RECT 23.18 135.09 157.32 136.8 ;
   RECT 23.18 136.8 157.32 138.51 ;
   RECT 23.18 138.51 157.32 140.22 ;
   RECT 23.18 140.22 157.32 141.93 ;
   RECT 23.18 141.93 157.32 143.64 ;
   RECT 23.18 143.64 157.32 145.35 ;
   RECT 23.18 145.35 157.32 147.06 ;
   RECT 23.18 147.06 157.32 148.77 ;
   RECT 23.18 148.77 157.32 150.48 ;
   RECT 23.18 150.48 157.32 152.19 ;
   RECT 23.18 152.19 157.32 153.9 ;
   RECT 23.18 153.9 157.32 155.61 ;
   RECT 23.18 155.61 157.32 157.32 ;
   RECT 23.18 157.32 157.32 159.03 ;
   RECT 23.18 159.03 157.32 160.74 ;
   RECT 23.18 160.74 157.32 162.45 ;
   RECT 23.18 162.45 157.32 164.16 ;
   RECT 23.18 164.16 157.32 165.87 ;
   RECT 23.18 165.87 157.32 167.58 ;
   RECT 23.18 167.58 157.32 169.29 ;
   RECT 23.18 169.29 157.32 171.0 ;
   RECT 23.18 171.0 157.32 172.71 ;
   RECT 23.18 172.71 157.32 174.42 ;
   RECT 23.18 174.42 157.32 176.13 ;
   RECT 23.18 176.13 157.32 177.84 ;
   RECT 0.0 177.84 157.32 179.55 ;
   RECT 0.0 179.55 157.32 181.26 ;
   RECT 0.0 181.26 157.32 182.97 ;
   RECT 0.0 182.97 157.32 184.68 ;
   RECT 0.0 184.68 157.32 186.39 ;
   RECT 0.0 186.39 157.32 188.1 ;
   RECT 0.0 188.1 157.32 189.81 ;
   RECT 0.0 189.81 157.32 191.52 ;
   RECT 0.0 191.52 157.32 193.23 ;
   RECT 0.0 193.23 157.32 194.94 ;
   RECT 0.0 194.94 157.32 196.65 ;
   RECT 0.0 196.65 157.32 198.36 ;
   RECT 0.0 198.36 157.32 200.07 ;
   RECT 0.0 200.07 157.32 201.78 ;
   RECT 0.0 201.78 157.32 203.49 ;
   RECT 0.0 203.49 157.32 205.2 ;
   RECT 0.0 205.2 157.32 206.91 ;
   RECT 23.18 206.91 157.32 208.62 ;
   RECT 23.18 208.62 157.32 210.33 ;
   RECT 23.18 210.33 157.32 212.04 ;
   RECT 23.18 212.04 157.32 213.75 ;
   RECT 23.18 213.75 157.32 215.46 ;
   RECT 23.18 215.46 157.32 217.17 ;
   RECT 23.18 217.17 157.32 218.88 ;
   RECT 23.18 218.88 157.32 220.59 ;
   RECT 23.18 220.59 157.32 222.3 ;
   RECT 23.18 222.3 157.32 224.01 ;
   RECT 23.18 224.01 157.32 225.72 ;
   RECT 23.18 225.72 157.32 227.43 ;
   RECT 23.18 227.43 157.32 229.14 ;
   RECT 23.18 229.14 157.32 230.85 ;
   RECT 23.18 230.85 157.32 232.56 ;
   RECT 23.18 232.56 157.32 234.27 ;
   RECT 23.18 234.27 157.32 235.98 ;
   RECT 23.18 235.98 157.32 237.69 ;
   RECT 23.18 237.69 157.32 239.4 ;
   RECT 23.18 239.4 157.32 241.11 ;
   RECT 23.18 241.11 157.32 242.82 ;
   RECT 23.18 242.82 157.32 244.53 ;
   RECT 23.18 244.53 157.32 246.24 ;
   RECT 23.18 246.24 157.32 247.95 ;
   RECT 23.18 247.95 157.32 249.66 ;
   RECT 23.18 249.66 157.32 251.37 ;
   RECT 23.18 251.37 157.32 253.08 ;
   RECT 23.18 253.08 157.32 254.79 ;
   RECT 23.18 254.79 157.32 256.5 ;
   RECT 23.18 256.5 157.32 258.21 ;
   RECT 23.18 258.21 157.32 259.92 ;
   RECT 23.18 259.92 157.32 261.63 ;
   RECT 23.18 261.63 157.32 263.34 ;
   RECT 23.18 263.34 157.32 265.05 ;
   RECT 23.18 265.05 157.32 266.76 ;
   RECT 23.18 266.76 157.32 268.47 ;
   RECT 23.18 268.47 157.32 270.18 ;
   RECT 23.18 270.18 157.32 271.89 ;
   RECT 23.18 271.89 157.32 273.6 ;
   RECT 23.18 273.6 157.32 275.31 ;
   RECT 23.18 275.31 157.32 277.02 ;
   RECT 23.18 277.02 157.32 278.73 ;
   RECT 23.18 278.73 157.32 280.44 ;
   RECT 23.18 280.44 157.32 282.15 ;
   RECT 23.18 282.15 157.32 283.86 ;
   RECT 23.18 283.86 157.32 285.57 ;
   RECT 23.18 285.57 157.32 287.28 ;
   RECT 23.18 287.28 157.32 288.99 ;
   RECT 23.18 288.99 157.32 290.7 ;
   RECT 23.18 290.7 157.32 292.41 ;
   RECT 23.18 292.41 157.32 294.12 ;
   RECT 23.18 294.12 157.32 295.83 ;
   RECT 23.18 295.83 157.32 297.54 ;
   RECT 23.18 297.54 157.32 299.25 ;
   RECT 23.18 299.25 157.32 300.96 ;
   RECT 23.18 300.96 157.32 302.67 ;
   RECT 23.18 302.67 157.32 304.38 ;
   RECT 23.18 304.38 157.32 306.09 ;
   RECT 23.18 306.09 157.32 307.8 ;
   RECT 23.18 307.8 157.32 309.51 ;
   RECT 23.18 309.51 157.32 311.22 ;
   RECT 23.18 311.22 157.32 312.93 ;
   RECT 23.18 312.93 157.32 314.64 ;
   RECT 23.18 314.64 157.32 316.35 ;
   RECT 23.18 316.35 157.32 318.06 ;
   RECT 23.18 318.06 157.32 319.77 ;
   RECT 23.18 319.77 157.32 321.48 ;
   RECT 23.18 321.48 157.32 323.19 ;
   RECT 23.18 323.19 157.32 324.9 ;
   RECT 23.18 324.9 157.32 326.61 ;
   RECT 23.18 326.61 157.32 328.32 ;
   RECT 23.18 328.32 157.32 330.03 ;
   RECT 23.18 330.03 157.32 331.74 ;
   RECT 23.18 331.74 157.32 333.45 ;
   RECT 23.18 333.45 157.32 335.16 ;
   RECT 23.18 335.16 157.32 336.87 ;
   RECT 23.18 336.87 157.32 338.58 ;
   RECT 23.18 338.58 157.32 340.29 ;
   RECT 23.18 340.29 157.32 342.0 ;
   RECT 23.18 342.0 157.32 343.71 ;
   RECT 23.18 343.71 157.32 345.42 ;
   RECT 23.18 345.42 157.32 347.13 ;
   RECT 23.18 347.13 157.32 348.84 ;
   RECT 23.18 348.84 157.32 350.55 ;
   RECT 23.18 350.55 157.32 352.26 ;
   RECT 23.18 352.26 157.32 353.97 ;
   RECT 23.18 353.97 157.32 355.68 ;
   RECT 23.18 355.68 157.32 357.39 ;
   RECT 23.18 357.39 157.32 359.1 ;
   RECT 23.18 359.1 157.32 360.81 ;
   RECT 23.18 360.81 157.32 362.52 ;
   RECT 23.18 362.52 157.32 364.23 ;
   RECT 23.18 364.23 157.32 365.94 ;
   RECT 23.18 365.94 157.32 367.65 ;
   RECT 23.18 367.65 157.32 369.36 ;
   RECT 23.18 369.36 157.32 371.07 ;
   RECT 23.18 371.07 157.32 372.78 ;
   RECT 23.18 372.78 157.32 374.49 ;
   RECT 23.18 374.49 157.32 376.2 ;
   RECT 23.18 376.2 157.32 377.91 ;
   RECT 23.18 377.91 157.32 379.62 ;
   RECT 23.18 379.62 157.32 381.33 ;
  LAYER via3 ;
   RECT 23.18 0.0 157.32 1.71 ;
   RECT 23.18 1.71 157.32 3.42 ;
   RECT 23.18 3.42 157.32 5.13 ;
   RECT 23.18 5.13 157.32 6.84 ;
   RECT 23.18 6.84 157.32 8.55 ;
   RECT 23.18 8.55 157.32 10.26 ;
   RECT 23.18 10.26 157.32 11.97 ;
   RECT 23.18 11.97 157.32 13.68 ;
   RECT 23.18 13.68 157.32 15.39 ;
   RECT 23.18 15.39 157.32 17.1 ;
   RECT 23.18 17.1 157.32 18.81 ;
   RECT 23.18 18.81 157.32 20.52 ;
   RECT 23.18 20.52 157.32 22.23 ;
   RECT 23.18 22.23 157.32 23.94 ;
   RECT 23.18 23.94 157.32 25.65 ;
   RECT 23.18 25.65 157.32 27.36 ;
   RECT 23.18 27.36 157.32 29.07 ;
   RECT 23.18 29.07 157.32 30.78 ;
   RECT 23.18 30.78 157.32 32.49 ;
   RECT 23.18 32.49 157.32 34.2 ;
   RECT 23.18 34.2 157.32 35.91 ;
   RECT 23.18 35.91 157.32 37.62 ;
   RECT 23.18 37.62 157.32 39.33 ;
   RECT 23.18 39.33 157.32 41.04 ;
   RECT 23.18 41.04 157.32 42.75 ;
   RECT 23.18 42.75 157.32 44.46 ;
   RECT 23.18 44.46 157.32 46.17 ;
   RECT 23.18 46.17 157.32 47.88 ;
   RECT 23.18 47.88 157.32 49.59 ;
   RECT 23.18 49.59 157.32 51.3 ;
   RECT 23.18 51.3 157.32 53.01 ;
   RECT 23.18 53.01 157.32 54.72 ;
   RECT 23.18 54.72 157.32 56.43 ;
   RECT 23.18 56.43 157.32 58.14 ;
   RECT 23.18 58.14 157.32 59.85 ;
   RECT 23.18 59.85 157.32 61.56 ;
   RECT 23.18 61.56 157.32 63.27 ;
   RECT 23.18 63.27 157.32 64.98 ;
   RECT 23.18 64.98 157.32 66.69 ;
   RECT 23.18 66.69 157.32 68.4 ;
   RECT 23.18 68.4 157.32 70.11 ;
   RECT 23.18 70.11 157.32 71.82 ;
   RECT 23.18 71.82 157.32 73.53 ;
   RECT 23.18 73.53 157.32 75.24 ;
   RECT 23.18 75.24 157.32 76.95 ;
   RECT 23.18 76.95 157.32 78.66 ;
   RECT 23.18 78.66 157.32 80.37 ;
   RECT 23.18 80.37 157.32 82.08 ;
   RECT 23.18 82.08 157.32 83.79 ;
   RECT 23.18 83.79 157.32 85.5 ;
   RECT 23.18 85.5 157.32 87.21 ;
   RECT 23.18 87.21 157.32 88.92 ;
   RECT 23.18 88.92 157.32 90.63 ;
   RECT 23.18 90.63 157.32 92.34 ;
   RECT 23.18 92.34 157.32 94.05 ;
   RECT 23.18 94.05 157.32 95.76 ;
   RECT 23.18 95.76 157.32 97.47 ;
   RECT 23.18 97.47 157.32 99.18 ;
   RECT 23.18 99.18 157.32 100.89 ;
   RECT 23.18 100.89 157.32 102.6 ;
   RECT 23.18 102.6 157.32 104.31 ;
   RECT 23.18 104.31 157.32 106.02 ;
   RECT 23.18 106.02 157.32 107.73 ;
   RECT 23.18 107.73 157.32 109.44 ;
   RECT 23.18 109.44 157.32 111.15 ;
   RECT 23.18 111.15 157.32 112.86 ;
   RECT 23.18 112.86 157.32 114.57 ;
   RECT 23.18 114.57 157.32 116.28 ;
   RECT 23.18 116.28 157.32 117.99 ;
   RECT 23.18 117.99 157.32 119.7 ;
   RECT 23.18 119.7 157.32 121.41 ;
   RECT 23.18 121.41 157.32 123.12 ;
   RECT 23.18 123.12 157.32 124.83 ;
   RECT 23.18 124.83 157.32 126.54 ;
   RECT 23.18 126.54 157.32 128.25 ;
   RECT 23.18 128.25 157.32 129.96 ;
   RECT 23.18 129.96 157.32 131.67 ;
   RECT 23.18 131.67 157.32 133.38 ;
   RECT 23.18 133.38 157.32 135.09 ;
   RECT 23.18 135.09 157.32 136.8 ;
   RECT 23.18 136.8 157.32 138.51 ;
   RECT 23.18 138.51 157.32 140.22 ;
   RECT 23.18 140.22 157.32 141.93 ;
   RECT 23.18 141.93 157.32 143.64 ;
   RECT 23.18 143.64 157.32 145.35 ;
   RECT 23.18 145.35 157.32 147.06 ;
   RECT 23.18 147.06 157.32 148.77 ;
   RECT 23.18 148.77 157.32 150.48 ;
   RECT 23.18 150.48 157.32 152.19 ;
   RECT 23.18 152.19 157.32 153.9 ;
   RECT 23.18 153.9 157.32 155.61 ;
   RECT 23.18 155.61 157.32 157.32 ;
   RECT 23.18 157.32 157.32 159.03 ;
   RECT 23.18 159.03 157.32 160.74 ;
   RECT 23.18 160.74 157.32 162.45 ;
   RECT 23.18 162.45 157.32 164.16 ;
   RECT 23.18 164.16 157.32 165.87 ;
   RECT 23.18 165.87 157.32 167.58 ;
   RECT 23.18 167.58 157.32 169.29 ;
   RECT 23.18 169.29 157.32 171.0 ;
   RECT 23.18 171.0 157.32 172.71 ;
   RECT 23.18 172.71 157.32 174.42 ;
   RECT 23.18 174.42 157.32 176.13 ;
   RECT 23.18 176.13 157.32 177.84 ;
   RECT 0.0 177.84 157.32 179.55 ;
   RECT 0.0 179.55 157.32 181.26 ;
   RECT 0.0 181.26 157.32 182.97 ;
   RECT 0.0 182.97 157.32 184.68 ;
   RECT 0.0 184.68 157.32 186.39 ;
   RECT 0.0 186.39 157.32 188.1 ;
   RECT 0.0 188.1 157.32 189.81 ;
   RECT 0.0 189.81 157.32 191.52 ;
   RECT 0.0 191.52 157.32 193.23 ;
   RECT 0.0 193.23 157.32 194.94 ;
   RECT 0.0 194.94 157.32 196.65 ;
   RECT 0.0 196.65 157.32 198.36 ;
   RECT 0.0 198.36 157.32 200.07 ;
   RECT 0.0 200.07 157.32 201.78 ;
   RECT 0.0 201.78 157.32 203.49 ;
   RECT 0.0 203.49 157.32 205.2 ;
   RECT 0.0 205.2 157.32 206.91 ;
   RECT 23.18 206.91 157.32 208.62 ;
   RECT 23.18 208.62 157.32 210.33 ;
   RECT 23.18 210.33 157.32 212.04 ;
   RECT 23.18 212.04 157.32 213.75 ;
   RECT 23.18 213.75 157.32 215.46 ;
   RECT 23.18 215.46 157.32 217.17 ;
   RECT 23.18 217.17 157.32 218.88 ;
   RECT 23.18 218.88 157.32 220.59 ;
   RECT 23.18 220.59 157.32 222.3 ;
   RECT 23.18 222.3 157.32 224.01 ;
   RECT 23.18 224.01 157.32 225.72 ;
   RECT 23.18 225.72 157.32 227.43 ;
   RECT 23.18 227.43 157.32 229.14 ;
   RECT 23.18 229.14 157.32 230.85 ;
   RECT 23.18 230.85 157.32 232.56 ;
   RECT 23.18 232.56 157.32 234.27 ;
   RECT 23.18 234.27 157.32 235.98 ;
   RECT 23.18 235.98 157.32 237.69 ;
   RECT 23.18 237.69 157.32 239.4 ;
   RECT 23.18 239.4 157.32 241.11 ;
   RECT 23.18 241.11 157.32 242.82 ;
   RECT 23.18 242.82 157.32 244.53 ;
   RECT 23.18 244.53 157.32 246.24 ;
   RECT 23.18 246.24 157.32 247.95 ;
   RECT 23.18 247.95 157.32 249.66 ;
   RECT 23.18 249.66 157.32 251.37 ;
   RECT 23.18 251.37 157.32 253.08 ;
   RECT 23.18 253.08 157.32 254.79 ;
   RECT 23.18 254.79 157.32 256.5 ;
   RECT 23.18 256.5 157.32 258.21 ;
   RECT 23.18 258.21 157.32 259.92 ;
   RECT 23.18 259.92 157.32 261.63 ;
   RECT 23.18 261.63 157.32 263.34 ;
   RECT 23.18 263.34 157.32 265.05 ;
   RECT 23.18 265.05 157.32 266.76 ;
   RECT 23.18 266.76 157.32 268.47 ;
   RECT 23.18 268.47 157.32 270.18 ;
   RECT 23.18 270.18 157.32 271.89 ;
   RECT 23.18 271.89 157.32 273.6 ;
   RECT 23.18 273.6 157.32 275.31 ;
   RECT 23.18 275.31 157.32 277.02 ;
   RECT 23.18 277.02 157.32 278.73 ;
   RECT 23.18 278.73 157.32 280.44 ;
   RECT 23.18 280.44 157.32 282.15 ;
   RECT 23.18 282.15 157.32 283.86 ;
   RECT 23.18 283.86 157.32 285.57 ;
   RECT 23.18 285.57 157.32 287.28 ;
   RECT 23.18 287.28 157.32 288.99 ;
   RECT 23.18 288.99 157.32 290.7 ;
   RECT 23.18 290.7 157.32 292.41 ;
   RECT 23.18 292.41 157.32 294.12 ;
   RECT 23.18 294.12 157.32 295.83 ;
   RECT 23.18 295.83 157.32 297.54 ;
   RECT 23.18 297.54 157.32 299.25 ;
   RECT 23.18 299.25 157.32 300.96 ;
   RECT 23.18 300.96 157.32 302.67 ;
   RECT 23.18 302.67 157.32 304.38 ;
   RECT 23.18 304.38 157.32 306.09 ;
   RECT 23.18 306.09 157.32 307.8 ;
   RECT 23.18 307.8 157.32 309.51 ;
   RECT 23.18 309.51 157.32 311.22 ;
   RECT 23.18 311.22 157.32 312.93 ;
   RECT 23.18 312.93 157.32 314.64 ;
   RECT 23.18 314.64 157.32 316.35 ;
   RECT 23.18 316.35 157.32 318.06 ;
   RECT 23.18 318.06 157.32 319.77 ;
   RECT 23.18 319.77 157.32 321.48 ;
   RECT 23.18 321.48 157.32 323.19 ;
   RECT 23.18 323.19 157.32 324.9 ;
   RECT 23.18 324.9 157.32 326.61 ;
   RECT 23.18 326.61 157.32 328.32 ;
   RECT 23.18 328.32 157.32 330.03 ;
   RECT 23.18 330.03 157.32 331.74 ;
   RECT 23.18 331.74 157.32 333.45 ;
   RECT 23.18 333.45 157.32 335.16 ;
   RECT 23.18 335.16 157.32 336.87 ;
   RECT 23.18 336.87 157.32 338.58 ;
   RECT 23.18 338.58 157.32 340.29 ;
   RECT 23.18 340.29 157.32 342.0 ;
   RECT 23.18 342.0 157.32 343.71 ;
   RECT 23.18 343.71 157.32 345.42 ;
   RECT 23.18 345.42 157.32 347.13 ;
   RECT 23.18 347.13 157.32 348.84 ;
   RECT 23.18 348.84 157.32 350.55 ;
   RECT 23.18 350.55 157.32 352.26 ;
   RECT 23.18 352.26 157.32 353.97 ;
   RECT 23.18 353.97 157.32 355.68 ;
   RECT 23.18 355.68 157.32 357.39 ;
   RECT 23.18 357.39 157.32 359.1 ;
   RECT 23.18 359.1 157.32 360.81 ;
   RECT 23.18 360.81 157.32 362.52 ;
   RECT 23.18 362.52 157.32 364.23 ;
   RECT 23.18 364.23 157.32 365.94 ;
   RECT 23.18 365.94 157.32 367.65 ;
   RECT 23.18 367.65 157.32 369.36 ;
   RECT 23.18 369.36 157.32 371.07 ;
   RECT 23.18 371.07 157.32 372.78 ;
   RECT 23.18 372.78 157.32 374.49 ;
   RECT 23.18 374.49 157.32 376.2 ;
   RECT 23.18 376.2 157.32 377.91 ;
   RECT 23.18 377.91 157.32 379.62 ;
   RECT 23.18 379.62 157.32 381.33 ;
  LAYER metal4 ;
   RECT 23.18 0.0 157.32 1.71 ;
   RECT 23.18 1.71 157.32 3.42 ;
   RECT 23.18 3.42 157.32 5.13 ;
   RECT 23.18 5.13 157.32 6.84 ;
   RECT 23.18 6.84 157.32 8.55 ;
   RECT 23.18 8.55 157.32 10.26 ;
   RECT 23.18 10.26 157.32 11.97 ;
   RECT 23.18 11.97 157.32 13.68 ;
   RECT 23.18 13.68 157.32 15.39 ;
   RECT 23.18 15.39 157.32 17.1 ;
   RECT 23.18 17.1 157.32 18.81 ;
   RECT 23.18 18.81 157.32 20.52 ;
   RECT 23.18 20.52 157.32 22.23 ;
   RECT 23.18 22.23 157.32 23.94 ;
   RECT 23.18 23.94 157.32 25.65 ;
   RECT 23.18 25.65 157.32 27.36 ;
   RECT 23.18 27.36 157.32 29.07 ;
   RECT 23.18 29.07 157.32 30.78 ;
   RECT 23.18 30.78 157.32 32.49 ;
   RECT 23.18 32.49 157.32 34.2 ;
   RECT 23.18 34.2 157.32 35.91 ;
   RECT 23.18 35.91 157.32 37.62 ;
   RECT 23.18 37.62 157.32 39.33 ;
   RECT 23.18 39.33 157.32 41.04 ;
   RECT 23.18 41.04 157.32 42.75 ;
   RECT 23.18 42.75 157.32 44.46 ;
   RECT 23.18 44.46 157.32 46.17 ;
   RECT 23.18 46.17 157.32 47.88 ;
   RECT 23.18 47.88 157.32 49.59 ;
   RECT 23.18 49.59 157.32 51.3 ;
   RECT 23.18 51.3 157.32 53.01 ;
   RECT 23.18 53.01 157.32 54.72 ;
   RECT 23.18 54.72 157.32 56.43 ;
   RECT 23.18 56.43 157.32 58.14 ;
   RECT 23.18 58.14 157.32 59.85 ;
   RECT 23.18 59.85 157.32 61.56 ;
   RECT 23.18 61.56 157.32 63.27 ;
   RECT 23.18 63.27 157.32 64.98 ;
   RECT 23.18 64.98 157.32 66.69 ;
   RECT 23.18 66.69 157.32 68.4 ;
   RECT 23.18 68.4 157.32 70.11 ;
   RECT 23.18 70.11 157.32 71.82 ;
   RECT 23.18 71.82 157.32 73.53 ;
   RECT 23.18 73.53 157.32 75.24 ;
   RECT 23.18 75.24 157.32 76.95 ;
   RECT 23.18 76.95 157.32 78.66 ;
   RECT 23.18 78.66 157.32 80.37 ;
   RECT 23.18 80.37 157.32 82.08 ;
   RECT 23.18 82.08 157.32 83.79 ;
   RECT 23.18 83.79 157.32 85.5 ;
   RECT 23.18 85.5 157.32 87.21 ;
   RECT 23.18 87.21 157.32 88.92 ;
   RECT 23.18 88.92 157.32 90.63 ;
   RECT 23.18 90.63 157.32 92.34 ;
   RECT 23.18 92.34 157.32 94.05 ;
   RECT 23.18 94.05 157.32 95.76 ;
   RECT 23.18 95.76 157.32 97.47 ;
   RECT 23.18 97.47 157.32 99.18 ;
   RECT 23.18 99.18 157.32 100.89 ;
   RECT 23.18 100.89 157.32 102.6 ;
   RECT 23.18 102.6 157.32 104.31 ;
   RECT 23.18 104.31 157.32 106.02 ;
   RECT 23.18 106.02 157.32 107.73 ;
   RECT 23.18 107.73 157.32 109.44 ;
   RECT 23.18 109.44 157.32 111.15 ;
   RECT 23.18 111.15 157.32 112.86 ;
   RECT 23.18 112.86 157.32 114.57 ;
   RECT 23.18 114.57 157.32 116.28 ;
   RECT 23.18 116.28 157.32 117.99 ;
   RECT 23.18 117.99 157.32 119.7 ;
   RECT 23.18 119.7 157.32 121.41 ;
   RECT 23.18 121.41 157.32 123.12 ;
   RECT 23.18 123.12 157.32 124.83 ;
   RECT 23.18 124.83 157.32 126.54 ;
   RECT 23.18 126.54 157.32 128.25 ;
   RECT 23.18 128.25 157.32 129.96 ;
   RECT 23.18 129.96 157.32 131.67 ;
   RECT 23.18 131.67 157.32 133.38 ;
   RECT 23.18 133.38 157.32 135.09 ;
   RECT 23.18 135.09 157.32 136.8 ;
   RECT 23.18 136.8 157.32 138.51 ;
   RECT 23.18 138.51 157.32 140.22 ;
   RECT 23.18 140.22 157.32 141.93 ;
   RECT 23.18 141.93 157.32 143.64 ;
   RECT 23.18 143.64 157.32 145.35 ;
   RECT 23.18 145.35 157.32 147.06 ;
   RECT 23.18 147.06 157.32 148.77 ;
   RECT 23.18 148.77 157.32 150.48 ;
   RECT 23.18 150.48 157.32 152.19 ;
   RECT 23.18 152.19 157.32 153.9 ;
   RECT 23.18 153.9 157.32 155.61 ;
   RECT 23.18 155.61 157.32 157.32 ;
   RECT 23.18 157.32 157.32 159.03 ;
   RECT 23.18 159.03 157.32 160.74 ;
   RECT 23.18 160.74 157.32 162.45 ;
   RECT 23.18 162.45 157.32 164.16 ;
   RECT 23.18 164.16 157.32 165.87 ;
   RECT 23.18 165.87 157.32 167.58 ;
   RECT 23.18 167.58 157.32 169.29 ;
   RECT 23.18 169.29 157.32 171.0 ;
   RECT 23.18 171.0 157.32 172.71 ;
   RECT 23.18 172.71 157.32 174.42 ;
   RECT 23.18 174.42 157.32 176.13 ;
   RECT 23.18 176.13 157.32 177.84 ;
   RECT 0.0 177.84 157.32 179.55 ;
   RECT 0.0 179.55 157.32 181.26 ;
   RECT 0.0 181.26 157.32 182.97 ;
   RECT 0.0 182.97 157.32 184.68 ;
   RECT 0.0 184.68 157.32 186.39 ;
   RECT 0.0 186.39 157.32 188.1 ;
   RECT 0.0 188.1 157.32 189.81 ;
   RECT 0.0 189.81 157.32 191.52 ;
   RECT 0.0 191.52 157.32 193.23 ;
   RECT 0.0 193.23 157.32 194.94 ;
   RECT 0.0 194.94 157.32 196.65 ;
   RECT 0.0 196.65 157.32 198.36 ;
   RECT 0.0 198.36 157.32 200.07 ;
   RECT 0.0 200.07 157.32 201.78 ;
   RECT 0.0 201.78 157.32 203.49 ;
   RECT 0.0 203.49 157.32 205.2 ;
   RECT 0.0 205.2 157.32 206.91 ;
   RECT 23.18 206.91 157.32 208.62 ;
   RECT 23.18 208.62 157.32 210.33 ;
   RECT 23.18 210.33 157.32 212.04 ;
   RECT 23.18 212.04 157.32 213.75 ;
   RECT 23.18 213.75 157.32 215.46 ;
   RECT 23.18 215.46 157.32 217.17 ;
   RECT 23.18 217.17 157.32 218.88 ;
   RECT 23.18 218.88 157.32 220.59 ;
   RECT 23.18 220.59 157.32 222.3 ;
   RECT 23.18 222.3 157.32 224.01 ;
   RECT 23.18 224.01 157.32 225.72 ;
   RECT 23.18 225.72 157.32 227.43 ;
   RECT 23.18 227.43 157.32 229.14 ;
   RECT 23.18 229.14 157.32 230.85 ;
   RECT 23.18 230.85 157.32 232.56 ;
   RECT 23.18 232.56 157.32 234.27 ;
   RECT 23.18 234.27 157.32 235.98 ;
   RECT 23.18 235.98 157.32 237.69 ;
   RECT 23.18 237.69 157.32 239.4 ;
   RECT 23.18 239.4 157.32 241.11 ;
   RECT 23.18 241.11 157.32 242.82 ;
   RECT 23.18 242.82 157.32 244.53 ;
   RECT 23.18 244.53 157.32 246.24 ;
   RECT 23.18 246.24 157.32 247.95 ;
   RECT 23.18 247.95 157.32 249.66 ;
   RECT 23.18 249.66 157.32 251.37 ;
   RECT 23.18 251.37 157.32 253.08 ;
   RECT 23.18 253.08 157.32 254.79 ;
   RECT 23.18 254.79 157.32 256.5 ;
   RECT 23.18 256.5 157.32 258.21 ;
   RECT 23.18 258.21 157.32 259.92 ;
   RECT 23.18 259.92 157.32 261.63 ;
   RECT 23.18 261.63 157.32 263.34 ;
   RECT 23.18 263.34 157.32 265.05 ;
   RECT 23.18 265.05 157.32 266.76 ;
   RECT 23.18 266.76 157.32 268.47 ;
   RECT 23.18 268.47 157.32 270.18 ;
   RECT 23.18 270.18 157.32 271.89 ;
   RECT 23.18 271.89 157.32 273.6 ;
   RECT 23.18 273.6 157.32 275.31 ;
   RECT 23.18 275.31 157.32 277.02 ;
   RECT 23.18 277.02 157.32 278.73 ;
   RECT 23.18 278.73 157.32 280.44 ;
   RECT 23.18 280.44 157.32 282.15 ;
   RECT 23.18 282.15 157.32 283.86 ;
   RECT 23.18 283.86 157.32 285.57 ;
   RECT 23.18 285.57 157.32 287.28 ;
   RECT 23.18 287.28 157.32 288.99 ;
   RECT 23.18 288.99 157.32 290.7 ;
   RECT 23.18 290.7 157.32 292.41 ;
   RECT 23.18 292.41 157.32 294.12 ;
   RECT 23.18 294.12 157.32 295.83 ;
   RECT 23.18 295.83 157.32 297.54 ;
   RECT 23.18 297.54 157.32 299.25 ;
   RECT 23.18 299.25 157.32 300.96 ;
   RECT 23.18 300.96 157.32 302.67 ;
   RECT 23.18 302.67 157.32 304.38 ;
   RECT 23.18 304.38 157.32 306.09 ;
   RECT 23.18 306.09 157.32 307.8 ;
   RECT 23.18 307.8 157.32 309.51 ;
   RECT 23.18 309.51 157.32 311.22 ;
   RECT 23.18 311.22 157.32 312.93 ;
   RECT 23.18 312.93 157.32 314.64 ;
   RECT 23.18 314.64 157.32 316.35 ;
   RECT 23.18 316.35 157.32 318.06 ;
   RECT 23.18 318.06 157.32 319.77 ;
   RECT 23.18 319.77 157.32 321.48 ;
   RECT 23.18 321.48 157.32 323.19 ;
   RECT 23.18 323.19 157.32 324.9 ;
   RECT 23.18 324.9 157.32 326.61 ;
   RECT 23.18 326.61 157.32 328.32 ;
   RECT 23.18 328.32 157.32 330.03 ;
   RECT 23.18 330.03 157.32 331.74 ;
   RECT 23.18 331.74 157.32 333.45 ;
   RECT 23.18 333.45 157.32 335.16 ;
   RECT 23.18 335.16 157.32 336.87 ;
   RECT 23.18 336.87 157.32 338.58 ;
   RECT 23.18 338.58 157.32 340.29 ;
   RECT 23.18 340.29 157.32 342.0 ;
   RECT 23.18 342.0 157.32 343.71 ;
   RECT 23.18 343.71 157.32 345.42 ;
   RECT 23.18 345.42 157.32 347.13 ;
   RECT 23.18 347.13 157.32 348.84 ;
   RECT 23.18 348.84 157.32 350.55 ;
   RECT 23.18 350.55 157.32 352.26 ;
   RECT 23.18 352.26 157.32 353.97 ;
   RECT 23.18 353.97 157.32 355.68 ;
   RECT 23.18 355.68 157.32 357.39 ;
   RECT 23.18 357.39 157.32 359.1 ;
   RECT 23.18 359.1 157.32 360.81 ;
   RECT 23.18 360.81 157.32 362.52 ;
   RECT 23.18 362.52 157.32 364.23 ;
   RECT 23.18 364.23 157.32 365.94 ;
   RECT 23.18 365.94 157.32 367.65 ;
   RECT 23.18 367.65 157.32 369.36 ;
   RECT 23.18 369.36 157.32 371.07 ;
   RECT 23.18 371.07 157.32 372.78 ;
   RECT 23.18 372.78 157.32 374.49 ;
   RECT 23.18 374.49 157.32 376.2 ;
   RECT 23.18 376.2 157.32 377.91 ;
   RECT 23.18 377.91 157.32 379.62 ;
   RECT 23.18 379.62 157.32 381.33 ;
 END
END block_414x2007_358

MACRO block_341x369_76
 CLASS BLOCK ;
 FOREIGN block_341x369_76 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 129.58 BY 70.11 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 20.235 126.445 20.805 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 26.695 126.445 27.265 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 6.935 3.325 7.505 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 9.215 3.325 9.785 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 10.735 3.325 11.305 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 13.015 3.325 13.585 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 13.395 4.085 13.965 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 13.775 3.325 14.345 ;
  END
 END o7
 PIN o8
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 15.295 3.325 15.865 ;
  END
 END o8
 PIN o9
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 16.055 3.325 16.625 ;
  END
 END o9
 PIN o10
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 64.315 29.735 64.885 30.305 ;
  END
 END o10
 PIN o11
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 12.635 4.085 13.205 ;
  END
 END o11
 PIN o12
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 19.855 3.325 20.425 ;
  END
 END o12
 PIN o13
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 20.615 3.325 21.185 ;
  END
 END o13
 PIN o14
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 21.375 3.325 21.945 ;
  END
 END o14
 PIN o15
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 22.135 3.325 22.705 ;
  END
 END o15
 PIN o16
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 64.315 28.975 64.885 29.545 ;
  END
 END o16
 PIN o17
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 18.335 3.325 18.905 ;
  END
 END o17
 PIN o18
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 25.935 3.325 26.505 ;
  END
 END o18
 PIN o19
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 26.695 3.325 27.265 ;
  END
 END o19
 PIN o20
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 27.455 3.325 28.025 ;
  END
 END o20
 PIN o21
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 28.975 3.325 29.545 ;
  END
 END o21
 PIN o22
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 65.075 29.735 65.645 30.305 ;
  END
 END o22
 PIN o23
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 25.175 3.325 25.745 ;
  END
 END o23
 PIN o24
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 32.015 3.325 32.585 ;
  END
 END o24
 PIN o25
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 33.535 3.325 34.105 ;
  END
 END o25
 PIN o26
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 34.295 3.325 34.865 ;
  END
 END o26
 PIN o27
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 35.055 3.325 35.625 ;
  END
 END o27
 PIN o28
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 64.315 35.055 64.885 35.625 ;
  END
 END o28
 PIN o29
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 31.255 3.325 31.825 ;
  END
 END o29
 PIN o30
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 38.095 126.445 38.665 ;
  END
 END o30
 PIN o31
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 38.855 126.445 39.425 ;
  END
 END o31
 PIN o32
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 39.615 126.445 40.185 ;
  END
 END o32
 PIN o33
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 21.755 126.445 22.325 ;
  END
 END o33
 PIN o34
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 31.255 126.445 31.825 ;
  END
 END o34
 PIN o35
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 32.015 126.445 32.585 ;
  END
 END o35
 PIN o36
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 33.535 126.445 34.105 ;
  END
 END o36
 PIN o37
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 30.495 126.445 31.065 ;
  END
 END o37
 PIN o38
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 28.975 126.445 29.545 ;
  END
 END o38
 PIN o39
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 41.135 3.325 41.705 ;
  END
 END o39
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 35.815 126.445 36.385 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 43.035 126.445 43.605 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 32.395 125.685 32.965 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 35.435 125.685 36.005 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 40.375 3.325 40.945 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 38.475 125.685 39.045 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 39.995 125.685 40.565 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 39.235 125.685 39.805 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 40.375 126.445 40.945 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 8.455 126.445 9.025 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 9.215 126.445 9.785 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 10.735 126.445 11.305 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 11.495 126.445 12.065 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 12.255 126.445 12.825 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 13.015 126.445 13.585 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 36.955 126.445 37.525 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 36.575 125.685 37.145 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 33.915 125.685 34.485 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 30.115 125.685 30.685 ;
  END
 END i18
 PIN i19
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 8.455 3.325 9.025 ;
  END
 END i19
 PIN i20
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 25.935 126.445 26.505 ;
  END
 END i20
 PIN i21
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 25.175 126.445 25.745 ;
  END
 END i21
 PIN i22
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 24.415 126.445 24.985 ;
  END
 END i22
 PIN i23
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 34.675 126.445 35.245 ;
  END
 END i23
 PIN i24
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 30.875 125.685 31.445 ;
  END
 END i24
 PIN i25
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 40.755 125.685 41.325 ;
  END
 END i25
 PIN i26
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 8.075 125.685 8.645 ;
  END
 END i26
 PIN i27
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 7.695 126.445 8.265 ;
  END
 END i27
 PIN i28
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 7.315 125.685 7.885 ;
  END
 END i28
 PIN i29
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 6.935 126.445 7.505 ;
  END
 END i29
 PIN i30
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 6.555 125.685 7.125 ;
  END
 END i30
 PIN i31
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 13.775 126.445 14.345 ;
  END
 END i31
 PIN i32
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 15.295 126.445 15.865 ;
  END
 END i32
 PIN i33
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 16.055 126.445 16.625 ;
  END
 END i33
 PIN i34
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 16.815 126.445 17.385 ;
  END
 END i34
 PIN i35
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 27.455 126.445 28.025 ;
  END
 END i35
 OBS
  LAYER metal1 ;
   RECT 0 0 129.58 70.11 ;
  LAYER via1 ;
   RECT 0 0 129.58 70.11 ;
  LAYER metal2 ;
   RECT 0 0 129.58 70.11 ;
  LAYER via2 ;
   RECT 0 0 129.58 70.11 ;
  LAYER metal3 ;
   RECT 0 0 129.58 70.11 ;
  LAYER via3 ;
   RECT 0 0 129.58 70.11 ;
  LAYER metal4 ;
   RECT 0 0 129.58 70.11 ;
 END
END block_341x369_76

MACRO block_737x1845_682
 CLASS BLOCK ;
 FOREIGN block_737x1845_682 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 280.06 BY 350.55 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 23.655 1.045 24.225 1.615 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 17.575 1.045 18.145 1.615 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 29.735 1.045 30.305 1.615 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 133.855 1.045 134.425 1.615 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 134.995 1.045 135.565 1.615 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 141.075 1.045 141.645 1.615 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 139.935 1.045 140.505 1.615 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 1.045 126.445 1.615 ;
  END
 END o7
 PIN o8
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 127.775 1.045 128.345 1.615 ;
  END
 END o8
 PIN o9
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 1.045 129.485 1.615 ;
  END
 END o9
 PIN o10
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 142.975 1.045 143.545 1.615 ;
  END
 END o10
 PIN o11
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 121.695 1.045 122.265 1.615 ;
  END
 END o11
 PIN o12
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 122.835 1.045 123.405 1.615 ;
  END
 END o12
 PIN o13
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 109.155 1.045 109.725 1.615 ;
  END
 END o13
 PIN o14
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 21.755 1.045 22.325 1.615 ;
  END
 END o14
 PIN o15
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.595 1.045 10.165 1.615 ;
  END
 END o15
 PIN o16
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 47.595 1.045 48.165 1.615 ;
  END
 END o16
 PIN o17
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 18.715 1.045 19.285 1.615 ;
  END
 END o17
 PIN o18
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 20.615 1.045 21.185 1.615 ;
  END
 END o18
 PIN o19
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 103.075 1.045 103.645 1.615 ;
  END
 END o19
 PIN o20
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 119.795 1.045 120.365 1.615 ;
  END
 END o20
 PIN o21
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 96.995 1.045 97.565 1.615 ;
  END
 END o21
 PIN o22
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 95.855 1.045 96.425 1.615 ;
  END
 END o22
 PIN o23
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 93.955 1.045 94.525 1.615 ;
  END
 END o23
 PIN o24
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 124.735 1.045 125.305 1.615 ;
  END
 END o24
 PIN o25
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.295 1.045 34.865 1.615 ;
  END
 END o25
 PIN o26
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 32.395 1.045 32.965 1.615 ;
  END
 END o26
 PIN o27
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 41.515 1.045 42.085 1.615 ;
  END
 END o27
 PIN o28
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 37.335 1.045 37.905 1.615 ;
  END
 END o28
 PIN o29
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 136.895 1.045 137.465 1.615 ;
  END
 END o29
 PIN o30
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 38.475 1.045 39.045 1.615 ;
  END
 END o30
 PIN o31
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 40.375 1.045 40.945 1.615 ;
  END
 END o31
 PIN o32
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 49.495 1.045 50.065 1.615 ;
  END
 END o32
 PIN o33
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 11.495 1.045 12.065 1.615 ;
  END
 END o33
 PIN o34
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 114.095 1.045 114.665 1.615 ;
  END
 END o34
 PIN o35
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.135 1.045 117.705 1.615 ;
  END
 END o35
 PIN o36
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 111.055 1.045 111.625 1.615 ;
  END
 END o36
 PIN o37
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 106.115 1.045 106.685 1.615 ;
  END
 END o37
 PIN o38
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 108.015 1.045 108.585 1.615 ;
  END
 END o38
 PIN o39
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 104.975 1.045 105.545 1.615 ;
  END
 END o39
 PIN o40
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 52.535 1.045 53.105 1.615 ;
  END
 END o40
 PIN o41
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.575 1.045 56.145 1.615 ;
  END
 END o41
 PIN o42
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 46.455 1.045 47.025 1.615 ;
  END
 END o42
 PIN o43
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 35.435 1.045 36.005 1.615 ;
  END
 END o43
 PIN o44
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 8.455 1.045 9.025 1.615 ;
  END
 END o44
 PIN o45
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 43.415 1.045 43.985 1.615 ;
  END
 END o45
 PIN o46
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 101.935 1.045 102.505 1.615 ;
  END
 END o46
 PIN o47
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 100.035 1.045 100.605 1.615 ;
  END
 END o47
 PIN o48
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 14.535 1.045 15.105 1.615 ;
  END
 END o48
 PIN o49
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 1.045 27.265 1.615 ;
  END
 END o49
 PIN o50
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 6.555 1.045 7.125 1.615 ;
  END
 END o50
 PIN o51
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 24.795 1.045 25.365 1.615 ;
  END
 END o51
 PIN o52
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 1.045 28.405 1.615 ;
  END
 END o52
 PIN o53
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 138.035 1.045 138.605 1.615 ;
  END
 END o53
 PIN o54
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 15.675 1.045 16.245 1.615 ;
  END
 END o54
 PIN o55
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 12.635 1.045 13.205 1.615 ;
  END
 END o55
 PIN o56
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 53.675 1.045 54.245 1.615 ;
  END
 END o56
 PIN o57
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 50.635 1.045 51.205 1.615 ;
  END
 END o57
 PIN o58
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 115.235 1.045 115.805 1.615 ;
  END
 END o58
 PIN o59
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 112.195 1.045 112.765 1.615 ;
  END
 END o59
 PIN o60
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 131.955 1.045 132.525 1.615 ;
  END
 END o60
 PIN o61
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 44.555 1.045 45.125 1.615 ;
  END
 END o61
 PIN o62
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 98.895 1.045 99.465 1.615 ;
  END
 END o62
 PIN o63
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.815 1.045 131.385 1.615 ;
  END
 END o63
 PIN o64
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 74.195 1.045 74.765 1.615 ;
  END
 END o64
 PIN o65
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 207.575 348.365 208.145 348.935 ;
  END
 END o65
 PIN o66
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.135 1.045 250.705 1.615 ;
  END
 END o66
 PIN o67
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 301.625 277.305 302.195 ;
  END
 END o67
 PIN o68
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 300.865 277.305 301.435 ;
  END
 END o68
 PIN o69
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 245.385 277.305 245.955 ;
  END
 END o69
 PIN o70
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 244.625 277.305 245.195 ;
  END
 END o70
 PIN o71
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 241.015 277.305 241.585 ;
  END
 END o71
 PIN o72
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 240.255 277.305 240.825 ;
  END
 END o72
 PIN o73
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 236.645 277.305 237.215 ;
  END
 END o73
 PIN o74
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 235.885 277.305 236.455 ;
  END
 END o74
 PIN o75
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 232.275 277.305 232.845 ;
  END
 END o75
 PIN o76
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 231.515 277.305 232.085 ;
  END
 END o76
 PIN o77
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 227.905 277.305 228.475 ;
  END
 END o77
 PIN o78
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 227.145 277.305 227.715 ;
  END
 END o78
 PIN o79
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 262.865 277.305 263.435 ;
  END
 END o79
 PIN o80
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 223.535 277.305 224.105 ;
  END
 END o80
 PIN o81
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 222.775 277.305 223.345 ;
  END
 END o81
 PIN o82
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 219.165 277.305 219.735 ;
  END
 END o82
 PIN o83
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 218.405 277.305 218.975 ;
  END
 END o83
 PIN o84
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 214.795 277.305 215.365 ;
  END
 END o84
 PIN o85
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 214.035 277.305 214.605 ;
  END
 END o85
 PIN o86
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 210.425 277.305 210.995 ;
  END
 END o86
 PIN o87
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 209.665 277.305 210.235 ;
  END
 END o87
 PIN o88
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 206.055 277.305 206.625 ;
  END
 END o88
 PIN o89
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 205.295 277.305 205.865 ;
  END
 END o89
 PIN o90
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 262.105 277.305 262.675 ;
  END
 END o90
 PIN o91
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 201.685 277.305 202.255 ;
  END
 END o91
 PIN o92
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 200.925 277.305 201.495 ;
  END
 END o92
 PIN o93
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 197.315 277.305 197.885 ;
  END
 END o93
 PIN o94
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 196.555 277.305 197.125 ;
  END
 END o94
 PIN o95
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 192.945 277.305 193.515 ;
  END
 END o95
 PIN o96
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 192.185 277.305 192.755 ;
  END
 END o96
 PIN o97
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 188.575 277.305 189.145 ;
  END
 END o97
 PIN o98
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 187.815 277.305 188.385 ;
  END
 END o98
 PIN o99
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 184.205 277.305 184.775 ;
  END
 END o99
 PIN o100
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 183.445 277.305 184.015 ;
  END
 END o100
 PIN o101
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 258.495 277.305 259.065 ;
  END
 END o101
 PIN o102
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 179.835 277.305 180.405 ;
  END
 END o102
 PIN o103
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 179.075 277.305 179.645 ;
  END
 END o103
 PIN o104
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 175.465 277.305 176.035 ;
  END
 END o104
 PIN o105
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 174.705 277.305 175.275 ;
  END
 END o105
 PIN o106
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 171.095 277.305 171.665 ;
  END
 END o106
 PIN o107
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 170.335 277.305 170.905 ;
  END
 END o107
 PIN o108
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 152.665 277.305 153.235 ;
  END
 END o108
 PIN o109
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 151.905 277.305 152.475 ;
  END
 END o109
 PIN o110
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 113.905 277.305 114.475 ;
  END
 END o110
 PIN o111
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 113.145 277.305 113.715 ;
  END
 END o111
 PIN o112
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 257.735 277.305 258.305 ;
  END
 END o112
 PIN o113
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 109.535 277.305 110.105 ;
  END
 END o113
 PIN o114
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 108.775 277.305 109.345 ;
  END
 END o114
 PIN o115
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 105.165 277.305 105.735 ;
  END
 END o115
 PIN o116
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 104.405 277.305 104.975 ;
  END
 END o116
 PIN o117
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 100.795 277.305 101.365 ;
  END
 END o117
 PIN o118
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 100.035 277.305 100.605 ;
  END
 END o118
 PIN o119
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 96.425 277.305 96.995 ;
  END
 END o119
 PIN o120
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 95.665 277.305 96.235 ;
  END
 END o120
 PIN o121
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 92.055 277.305 92.625 ;
  END
 END o121
 PIN o122
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 91.295 277.305 91.865 ;
  END
 END o122
 PIN o123
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 254.125 277.305 254.695 ;
  END
 END o123
 PIN o124
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 87.685 277.305 88.255 ;
  END
 END o124
 PIN o125
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 86.925 277.305 87.495 ;
  END
 END o125
 PIN o126
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 83.315 277.305 83.885 ;
  END
 END o126
 PIN o127
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 82.555 277.305 83.125 ;
  END
 END o127
 PIN o128
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 78.945 277.305 79.515 ;
  END
 END o128
 PIN o129
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 78.185 277.305 78.755 ;
  END
 END o129
 PIN o130
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 74.575 277.305 75.145 ;
  END
 END o130
 PIN o131
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 73.815 277.305 74.385 ;
  END
 END o131
 PIN o132
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 70.205 277.305 70.775 ;
  END
 END o132
 PIN o133
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 69.445 277.305 70.015 ;
  END
 END o133
 PIN o134
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 253.365 277.305 253.935 ;
  END
 END o134
 PIN o135
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 65.835 277.305 66.405 ;
  END
 END o135
 PIN o136
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 65.075 277.305 65.645 ;
  END
 END o136
 PIN o137
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 61.465 277.305 62.035 ;
  END
 END o137
 PIN o138
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 60.705 277.305 61.275 ;
  END
 END o138
 PIN o139
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 57.095 277.305 57.665 ;
  END
 END o139
 PIN o140
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 56.335 277.305 56.905 ;
  END
 END o140
 PIN o141
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 52.725 277.305 53.295 ;
  END
 END o141
 PIN o142
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 51.965 277.305 52.535 ;
  END
 END o142
 PIN o143
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 48.355 277.305 48.925 ;
  END
 END o143
 PIN o144
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 47.595 277.305 48.165 ;
  END
 END o144
 PIN o145
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 249.755 277.305 250.325 ;
  END
 END o145
 PIN o146
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 43.985 277.305 44.555 ;
  END
 END o146
 PIN o147
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 43.225 277.305 43.795 ;
  END
 END o147
 PIN o148
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 39.615 277.305 40.185 ;
  END
 END o148
 PIN o149
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 38.855 277.305 39.425 ;
  END
 END o149
 PIN o150
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 35.245 277.305 35.815 ;
  END
 END o150
 PIN o151
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 34.485 277.305 35.055 ;
  END
 END o151
 PIN o152
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 30.875 277.305 31.445 ;
  END
 END o152
 PIN o153
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 30.115 277.305 30.685 ;
  END
 END o153
 PIN o154
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 26.505 277.305 27.075 ;
  END
 END o154
 PIN o155
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 25.745 277.305 26.315 ;
  END
 END o155
 PIN o156
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 248.995 277.305 249.565 ;
  END
 END o156
 PIN o157
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 22.135 277.305 22.705 ;
  END
 END o157
 PIN o158
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 21.375 277.305 21.945 ;
  END
 END o158
 PIN o159
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 302.195 251.465 302.765 ;
  END
 END o159
 PIN o160
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 299.915 251.465 300.485 ;
  END
 END o160
 PIN o161
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 245.575 251.465 246.145 ;
  END
 END o161
 PIN o162
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 244.245 251.465 244.815 ;
  END
 END o162
 PIN o163
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 241.205 251.465 241.775 ;
  END
 END o163
 PIN o164
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 239.875 251.465 240.445 ;
  END
 END o164
 PIN o165
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 236.835 251.465 237.405 ;
  END
 END o165
 PIN o166
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 235.505 251.465 236.075 ;
  END
 END o166
 PIN o167
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 232.465 251.465 233.035 ;
  END
 END o167
 PIN o168
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 231.135 251.465 231.705 ;
  END
 END o168
 PIN o169
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 228.095 251.465 228.665 ;
  END
 END o169
 PIN o170
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 226.765 251.465 227.335 ;
  END
 END o170
 PIN o171
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 263.055 251.465 263.625 ;
  END
 END o171
 PIN o172
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 223.725 251.465 224.295 ;
  END
 END o172
 PIN o173
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 222.395 251.465 222.965 ;
  END
 END o173
 PIN o174
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 219.355 251.465 219.925 ;
  END
 END o174
 PIN o175
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 218.025 251.465 218.595 ;
  END
 END o175
 PIN o176
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 214.985 251.465 215.555 ;
  END
 END o176
 PIN o177
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 213.655 251.465 214.225 ;
  END
 END o177
 PIN o178
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 210.615 251.465 211.185 ;
  END
 END o178
 PIN o179
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 209.285 251.465 209.855 ;
  END
 END o179
 PIN o180
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 206.245 251.465 206.815 ;
  END
 END o180
 PIN o181
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 204.915 251.465 205.485 ;
  END
 END o181
 PIN o182
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 261.725 251.465 262.295 ;
  END
 END o182
 PIN o183
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 201.875 251.465 202.445 ;
  END
 END o183
 PIN o184
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 200.545 251.465 201.115 ;
  END
 END o184
 PIN o185
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 197.505 251.465 198.075 ;
  END
 END o185
 PIN o186
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 196.175 251.465 196.745 ;
  END
 END o186
 PIN o187
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 193.135 251.465 193.705 ;
  END
 END o187
 PIN o188
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 191.805 251.465 192.375 ;
  END
 END o188
 PIN o189
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 188.765 251.465 189.335 ;
  END
 END o189
 PIN o190
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 187.435 251.465 188.005 ;
  END
 END o190
 PIN o191
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 184.395 251.465 184.965 ;
  END
 END o191
 PIN o192
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 183.065 251.465 183.635 ;
  END
 END o192
 PIN o193
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 258.685 251.465 259.255 ;
  END
 END o193
 PIN o194
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 180.025 251.465 180.595 ;
  END
 END o194
 PIN o195
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 178.695 251.465 179.265 ;
  END
 END o195
 PIN o196
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 175.655 251.465 176.225 ;
  END
 END o196
 PIN o197
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 174.325 251.465 174.895 ;
  END
 END o197
 PIN o198
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 171.285 251.465 171.855 ;
  END
 END o198
 PIN o199
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 169.955 251.465 170.525 ;
  END
 END o199
 PIN o200
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 153.235 251.465 153.805 ;
  END
 END o200
 PIN o201
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 150.955 251.465 151.525 ;
  END
 END o201
 PIN o202
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 114.095 251.465 114.665 ;
  END
 END o202
 PIN o203
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 112.765 251.465 113.335 ;
  END
 END o203
 PIN o204
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 257.355 251.465 257.925 ;
  END
 END o204
 PIN o205
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 109.725 251.465 110.295 ;
  END
 END o205
 PIN o206
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 108.395 251.465 108.965 ;
  END
 END o206
 PIN o207
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 105.355 251.465 105.925 ;
  END
 END o207
 PIN o208
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 104.025 251.465 104.595 ;
  END
 END o208
 PIN o209
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 100.985 251.465 101.555 ;
  END
 END o209
 PIN o210
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 99.655 251.465 100.225 ;
  END
 END o210
 PIN o211
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 96.615 251.465 97.185 ;
  END
 END o211
 PIN o212
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 95.285 251.465 95.855 ;
  END
 END o212
 PIN o213
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 92.245 251.465 92.815 ;
  END
 END o213
 PIN o214
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 90.915 251.465 91.485 ;
  END
 END o214
 PIN o215
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 254.315 251.465 254.885 ;
  END
 END o215
 PIN o216
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 87.875 251.465 88.445 ;
  END
 END o216
 PIN o217
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 86.545 251.465 87.115 ;
  END
 END o217
 PIN o218
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 83.505 251.465 84.075 ;
  END
 END o218
 PIN o219
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 82.175 251.465 82.745 ;
  END
 END o219
 PIN o220
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 79.135 251.465 79.705 ;
  END
 END o220
 PIN o221
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 77.805 251.465 78.375 ;
  END
 END o221
 PIN o222
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 74.765 251.465 75.335 ;
  END
 END o222
 PIN o223
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 73.435 251.465 74.005 ;
  END
 END o223
 PIN o224
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 70.395 251.465 70.965 ;
  END
 END o224
 PIN o225
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 69.065 251.465 69.635 ;
  END
 END o225
 PIN o226
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 252.985 251.465 253.555 ;
  END
 END o226
 PIN o227
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 66.025 251.465 66.595 ;
  END
 END o227
 PIN o228
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 64.695 251.465 65.265 ;
  END
 END o228
 PIN o229
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 61.655 251.465 62.225 ;
  END
 END o229
 PIN o230
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 60.325 251.465 60.895 ;
  END
 END o230
 PIN o231
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 57.285 251.465 57.855 ;
  END
 END o231
 PIN o232
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 55.955 251.465 56.525 ;
  END
 END o232
 PIN o233
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 52.915 251.465 53.485 ;
  END
 END o233
 PIN o234
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 51.585 251.465 52.155 ;
  END
 END o234
 PIN o235
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 48.545 251.465 49.115 ;
  END
 END o235
 PIN o236
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 47.215 251.465 47.785 ;
  END
 END o236
 PIN o237
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 249.945 251.465 250.515 ;
  END
 END o237
 PIN o238
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 44.175 251.465 44.745 ;
  END
 END o238
 PIN o239
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 42.845 251.465 43.415 ;
  END
 END o239
 PIN o240
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 39.805 251.465 40.375 ;
  END
 END o240
 PIN o241
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 38.475 251.465 39.045 ;
  END
 END o241
 PIN o242
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 35.435 251.465 36.005 ;
  END
 END o242
 PIN o243
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 34.105 251.465 34.675 ;
  END
 END o243
 PIN o244
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 31.065 251.465 31.635 ;
  END
 END o244
 PIN o245
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 29.735 251.465 30.305 ;
  END
 END o245
 PIN o246
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 26.695 251.465 27.265 ;
  END
 END o246
 PIN o247
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 25.365 251.465 25.935 ;
  END
 END o247
 PIN o248
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 248.615 251.465 249.185 ;
  END
 END o248
 PIN o249
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 22.325 251.465 22.895 ;
  END
 END o249
 PIN o250
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 20.995 251.465 21.565 ;
  END
 END o250
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 235.315 348.365 235.885 348.935 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 223.155 348.365 223.725 348.935 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 224.675 348.365 225.245 348.935 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 236.075 348.365 236.645 348.935 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 223.915 348.365 224.485 348.935 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 237.215 348.365 237.785 348.935 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 248.235 269.705 248.805 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 20.615 269.705 21.185 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 22.705 269.705 23.275 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 250.325 269.705 250.895 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 24.985 269.705 25.555 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 27.075 269.705 27.645 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 29.355 269.705 29.925 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 31.445 269.705 32.015 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 33.725 269.705 34.295 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 35.815 269.705 36.385 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 38.095 269.705 38.665 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 40.185 269.705 40.755 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 42.465 269.705 43.035 ;
  END
 END i18
 PIN i19
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 44.555 269.705 45.125 ;
  END
 END i19
 PIN i20
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 252.605 269.705 253.175 ;
  END
 END i20
 PIN i21
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 46.835 269.705 47.405 ;
  END
 END i21
 PIN i22
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 48.925 269.705 49.495 ;
  END
 END i22
 PIN i23
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 51.205 269.705 51.775 ;
  END
 END i23
 PIN i24
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 53.295 269.705 53.865 ;
  END
 END i24
 PIN i25
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 55.575 269.705 56.145 ;
  END
 END i25
 PIN i26
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 57.665 269.705 58.235 ;
  END
 END i26
 PIN i27
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 59.945 269.705 60.515 ;
  END
 END i27
 PIN i28
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 62.035 269.705 62.605 ;
  END
 END i28
 PIN i29
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 64.315 269.705 64.885 ;
  END
 END i29
 PIN i30
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 66.405 269.705 66.975 ;
  END
 END i30
 PIN i31
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 254.695 269.705 255.265 ;
  END
 END i31
 PIN i32
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 70.775 269.705 71.345 ;
  END
 END i32
 PIN i33
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 73.055 269.705 73.625 ;
  END
 END i33
 PIN i34
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 75.145 269.705 75.715 ;
  END
 END i34
 PIN i35
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 77.425 269.705 77.995 ;
  END
 END i35
 PIN i36
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 79.515 269.705 80.085 ;
  END
 END i36
 PIN i37
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 81.795 269.705 82.365 ;
  END
 END i37
 PIN i38
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 83.885 269.705 84.455 ;
  END
 END i38
 PIN i39
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 86.165 269.705 86.735 ;
  END
 END i39
 PIN i40
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 88.255 269.705 88.825 ;
  END
 END i40
 PIN i41
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 256.975 269.705 257.545 ;
  END
 END i41
 PIN i42
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 90.535 269.705 91.105 ;
  END
 END i42
 PIN i43
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 92.625 269.705 93.195 ;
  END
 END i43
 PIN i44
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 94.905 269.705 95.475 ;
  END
 END i44
 PIN i45
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 96.995 269.705 97.565 ;
  END
 END i45
 PIN i46
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 99.275 269.705 99.845 ;
  END
 END i46
 PIN i47
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 101.365 269.705 101.935 ;
  END
 END i47
 PIN i48
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 103.645 269.705 104.215 ;
  END
 END i48
 PIN i49
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 105.735 269.705 106.305 ;
  END
 END i49
 PIN i50
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 108.015 269.705 108.585 ;
  END
 END i50
 PIN i51
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 110.105 269.705 110.675 ;
  END
 END i51
 PIN i52
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 259.065 269.705 259.635 ;
  END
 END i52
 PIN i53
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 112.385 269.705 112.955 ;
  END
 END i53
 PIN i54
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 114.475 269.705 115.045 ;
  END
 END i54
 PIN i55
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 150.955 269.705 151.525 ;
  END
 END i55
 PIN i56
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 153.045 269.705 153.615 ;
  END
 END i56
 PIN i57
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 171.665 269.705 172.235 ;
  END
 END i57
 PIN i58
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 176.035 269.705 176.605 ;
  END
 END i58
 PIN i59
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 180.405 269.705 180.975 ;
  END
 END i59
 PIN i60
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 261.345 269.705 261.915 ;
  END
 END i60
 PIN i61
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 182.685 269.705 183.255 ;
  END
 END i61
 PIN i62
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 184.775 269.705 185.345 ;
  END
 END i62
 PIN i63
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 187.055 269.705 187.625 ;
  END
 END i63
 PIN i64
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 189.145 269.705 189.715 ;
  END
 END i64
 PIN i65
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 191.425 269.705 191.995 ;
  END
 END i65
 PIN i66
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 193.515 269.705 194.085 ;
  END
 END i66
 PIN i67
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 195.795 269.705 196.365 ;
  END
 END i67
 PIN i68
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 197.885 269.705 198.455 ;
  END
 END i68
 PIN i69
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 200.165 269.705 200.735 ;
  END
 END i69
 PIN i70
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 202.255 269.705 202.825 ;
  END
 END i70
 PIN i71
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 263.435 269.705 264.005 ;
  END
 END i71
 PIN i72
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 204.535 269.705 205.105 ;
  END
 END i72
 PIN i73
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 206.625 269.705 207.195 ;
  END
 END i73
 PIN i74
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 208.905 269.705 209.475 ;
  END
 END i74
 PIN i75
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 210.995 269.705 211.565 ;
  END
 END i75
 PIN i76
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 213.275 269.705 213.845 ;
  END
 END i76
 PIN i77
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 215.365 269.705 215.935 ;
  END
 END i77
 PIN i78
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 217.645 269.705 218.215 ;
  END
 END i78
 PIN i79
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 219.735 269.705 220.305 ;
  END
 END i79
 PIN i80
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 222.015 269.705 222.585 ;
  END
 END i80
 PIN i81
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 224.105 269.705 224.675 ;
  END
 END i81
 PIN i82
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 299.915 269.705 300.485 ;
  END
 END i82
 PIN i83
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 226.385 269.705 226.955 ;
  END
 END i83
 PIN i84
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 228.475 269.705 229.045 ;
  END
 END i84
 PIN i85
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 230.755 269.705 231.325 ;
  END
 END i85
 PIN i86
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 232.845 269.705 233.415 ;
  END
 END i86
 PIN i87
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 235.125 269.705 235.695 ;
  END
 END i87
 PIN i88
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 237.215 269.705 237.785 ;
  END
 END i88
 PIN i89
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 239.495 269.705 240.065 ;
  END
 END i89
 PIN i90
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 241.585 269.705 242.155 ;
  END
 END i90
 PIN i91
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 243.865 269.705 244.435 ;
  END
 END i91
 PIN i92
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 245.955 269.705 246.525 ;
  END
 END i92
 PIN i93
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 302.005 269.705 302.575 ;
  END
 END i93
 PIN i94
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 173.945 269.705 174.515 ;
  END
 END i94
 PIN i95
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 169.575 269.705 170.145 ;
  END
 END i95
 PIN i96
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 178.315 269.705 178.885 ;
  END
 END i96
 PIN i97
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 68.685 269.705 69.255 ;
  END
 END i97
 PIN i98
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 220.115 348.365 220.685 348.935 ;
  END
 END i98
 PIN i99
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.775 348.365 242.345 348.935 ;
  END
 END i99
 PIN i100
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 243.675 348.365 244.245 348.935 ;
  END
 END i100
 PIN i101
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 218.595 348.365 219.165 348.935 ;
  END
 END i101
 PIN i102
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 239.875 348.365 240.445 348.935 ;
  END
 END i102
 PIN i103
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 245.195 348.365 245.765 348.935 ;
  END
 END i103
 PIN i104
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 209.475 348.365 210.045 348.935 ;
  END
 END i104
 PIN i105
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 208.335 348.365 208.905 348.935 ;
  END
 END i105
 PIN i106
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.635 348.365 241.205 348.935 ;
  END
 END i106
 PIN i107
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 217.455 348.365 218.025 348.935 ;
  END
 END i107
 PIN i108
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 219.355 348.365 219.925 348.935 ;
  END
 END i108
 PIN i109
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 244.435 348.365 245.005 348.935 ;
  END
 END i109
 PIN i110
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 242.535 348.365 243.105 348.935 ;
  END
 END i110
 PIN i111
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 302.005 276.545 302.575 ;
  END
 END i111
 PIN i112
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 300.295 276.545 300.865 ;
  END
 END i112
 PIN i113
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 245.765 276.545 246.335 ;
  END
 END i113
 PIN i114
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 244.055 276.545 244.625 ;
  END
 END i114
 PIN i115
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 241.395 276.545 241.965 ;
  END
 END i115
 PIN i116
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 239.685 276.545 240.255 ;
  END
 END i116
 PIN i117
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 237.025 276.545 237.595 ;
  END
 END i117
 PIN i118
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 235.315 276.545 235.885 ;
  END
 END i118
 PIN i119
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 232.655 276.545 233.225 ;
  END
 END i119
 PIN i120
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 230.945 276.545 231.515 ;
  END
 END i120
 PIN i121
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 228.285 276.545 228.855 ;
  END
 END i121
 PIN i122
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 226.575 276.545 227.145 ;
  END
 END i122
 PIN i123
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 263.245 276.545 263.815 ;
  END
 END i123
 PIN i124
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 223.915 276.545 224.485 ;
  END
 END i124
 PIN i125
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 222.205 276.545 222.775 ;
  END
 END i125
 PIN i126
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 219.545 276.545 220.115 ;
  END
 END i126
 PIN i127
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 217.835 276.545 218.405 ;
  END
 END i127
 PIN i128
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 215.175 276.545 215.745 ;
  END
 END i128
 PIN i129
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 213.465 276.545 214.035 ;
  END
 END i129
 PIN i130
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 210.805 276.545 211.375 ;
  END
 END i130
 PIN i131
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 209.095 276.545 209.665 ;
  END
 END i131
 PIN i132
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 206.435 276.545 207.005 ;
  END
 END i132
 PIN i133
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 204.725 276.545 205.295 ;
  END
 END i133
 PIN i134
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 261.535 276.545 262.105 ;
  END
 END i134
 PIN i135
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 202.065 276.545 202.635 ;
  END
 END i135
 PIN i136
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 200.355 276.545 200.925 ;
  END
 END i136
 PIN i137
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 197.695 276.545 198.265 ;
  END
 END i137
 PIN i138
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 195.985 276.545 196.555 ;
  END
 END i138
 PIN i139
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 193.325 276.545 193.895 ;
  END
 END i139
 PIN i140
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 191.615 276.545 192.185 ;
  END
 END i140
 PIN i141
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 188.955 276.545 189.525 ;
  END
 END i141
 PIN i142
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 187.245 276.545 187.815 ;
  END
 END i142
 PIN i143
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 184.585 276.545 185.155 ;
  END
 END i143
 PIN i144
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 182.875 276.545 183.445 ;
  END
 END i144
 PIN i145
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 258.875 276.545 259.445 ;
  END
 END i145
 PIN i146
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 180.215 276.545 180.785 ;
  END
 END i146
 PIN i147
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 178.505 276.545 179.075 ;
  END
 END i147
 PIN i148
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 175.845 276.545 176.415 ;
  END
 END i148
 PIN i149
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 174.135 276.545 174.705 ;
  END
 END i149
 PIN i150
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 171.475 276.545 172.045 ;
  END
 END i150
 PIN i151
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 169.765 276.545 170.335 ;
  END
 END i151
 PIN i152
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 153.235 276.545 153.805 ;
  END
 END i152
 PIN i153
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 151.525 276.545 152.095 ;
  END
 END i153
 PIN i154
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 114.285 276.545 114.855 ;
  END
 END i154
 PIN i155
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 112.575 276.545 113.145 ;
  END
 END i155
 PIN i156
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 257.165 276.545 257.735 ;
  END
 END i156
 PIN i157
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 109.915 276.545 110.485 ;
  END
 END i157
 PIN i158
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 108.205 276.545 108.775 ;
  END
 END i158
 PIN i159
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 105.545 276.545 106.115 ;
  END
 END i159
 PIN i160
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 103.835 276.545 104.405 ;
  END
 END i160
 PIN i161
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 101.175 276.545 101.745 ;
  END
 END i161
 PIN i162
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 99.465 276.545 100.035 ;
  END
 END i162
 PIN i163
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 96.805 276.545 97.375 ;
  END
 END i163
 PIN i164
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 95.095 276.545 95.665 ;
  END
 END i164
 PIN i165
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 92.435 276.545 93.005 ;
  END
 END i165
 PIN i166
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 90.725 276.545 91.295 ;
  END
 END i166
 PIN i167
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 254.505 276.545 255.075 ;
  END
 END i167
 PIN i168
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 88.065 276.545 88.635 ;
  END
 END i168
 PIN i169
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 86.355 276.545 86.925 ;
  END
 END i169
 PIN i170
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 83.695 276.545 84.265 ;
  END
 END i170
 PIN i171
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 81.985 276.545 82.555 ;
  END
 END i171
 PIN i172
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 79.325 276.545 79.895 ;
  END
 END i172
 PIN i173
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 77.615 276.545 78.185 ;
  END
 END i173
 PIN i174
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 74.955 276.545 75.525 ;
  END
 END i174
 PIN i175
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 73.245 276.545 73.815 ;
  END
 END i175
 PIN i176
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 70.585 276.545 71.155 ;
  END
 END i176
 PIN i177
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 68.875 276.545 69.445 ;
  END
 END i177
 PIN i178
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 252.795 276.545 253.365 ;
  END
 END i178
 PIN i179
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 66.215 276.545 66.785 ;
  END
 END i179
 PIN i180
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 64.505 276.545 65.075 ;
  END
 END i180
 PIN i181
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 61.845 276.545 62.415 ;
  END
 END i181
 PIN i182
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 60.135 276.545 60.705 ;
  END
 END i182
 PIN i183
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 57.475 276.545 58.045 ;
  END
 END i183
 PIN i184
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 55.765 276.545 56.335 ;
  END
 END i184
 PIN i185
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 53.105 276.545 53.675 ;
  END
 END i185
 PIN i186
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 51.395 276.545 51.965 ;
  END
 END i186
 PIN i187
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 48.735 276.545 49.305 ;
  END
 END i187
 PIN i188
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 47.025 276.545 47.595 ;
  END
 END i188
 PIN i189
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 250.135 276.545 250.705 ;
  END
 END i189
 PIN i190
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 44.365 276.545 44.935 ;
  END
 END i190
 PIN i191
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 42.655 276.545 43.225 ;
  END
 END i191
 PIN i192
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 39.995 276.545 40.565 ;
  END
 END i192
 PIN i193
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 38.285 276.545 38.855 ;
  END
 END i193
 PIN i194
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 35.625 276.545 36.195 ;
  END
 END i194
 PIN i195
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 33.915 276.545 34.485 ;
  END
 END i195
 PIN i196
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 31.255 276.545 31.825 ;
  END
 END i196
 PIN i197
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 29.545 276.545 30.115 ;
  END
 END i197
 PIN i198
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 26.885 276.545 27.455 ;
  END
 END i198
 PIN i199
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 25.175 276.545 25.745 ;
  END
 END i199
 PIN i200
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 248.425 276.545 248.995 ;
  END
 END i200
 PIN i201
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 22.515 276.545 23.085 ;
  END
 END i201
 PIN i202
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 20.805 276.545 21.375 ;
  END
 END i202
 PIN i203
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 302.575 277.305 303.145 ;
  END
 END i203
 PIN i204
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 299.915 277.305 300.485 ;
  END
 END i204
 PIN i205
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 246.335 277.305 246.905 ;
  END
 END i205
 PIN i206
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 243.675 277.305 244.245 ;
  END
 END i206
 PIN i207
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 241.965 277.305 242.535 ;
  END
 END i207
 PIN i208
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 239.305 277.305 239.875 ;
  END
 END i208
 PIN i209
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 237.595 277.305 238.165 ;
  END
 END i209
 PIN i210
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 234.935 277.305 235.505 ;
  END
 END i210
 PIN i211
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 233.225 277.305 233.795 ;
  END
 END i211
 PIN i212
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 230.565 277.305 231.135 ;
  END
 END i212
 PIN i213
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 228.855 277.305 229.425 ;
  END
 END i213
 PIN i214
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 226.195 277.305 226.765 ;
  END
 END i214
 PIN i215
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 263.815 277.305 264.385 ;
  END
 END i215
 PIN i216
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 224.485 277.305 225.055 ;
  END
 END i216
 PIN i217
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 221.825 277.305 222.395 ;
  END
 END i217
 PIN i218
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 220.115 277.305 220.685 ;
  END
 END i218
 PIN i219
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 217.455 277.305 218.025 ;
  END
 END i219
 PIN i220
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 215.745 277.305 216.315 ;
  END
 END i220
 PIN i221
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 213.085 277.305 213.655 ;
  END
 END i221
 PIN i222
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 211.375 277.305 211.945 ;
  END
 END i222
 PIN i223
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 208.715 277.305 209.285 ;
  END
 END i223
 PIN i224
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 207.005 277.305 207.575 ;
  END
 END i224
 PIN i225
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 204.345 277.305 204.915 ;
  END
 END i225
 PIN i226
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 261.155 277.305 261.725 ;
  END
 END i226
 PIN i227
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 202.635 277.305 203.205 ;
  END
 END i227
 PIN i228
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 199.975 277.305 200.545 ;
  END
 END i228
 PIN i229
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 198.265 277.305 198.835 ;
  END
 END i229
 PIN i230
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 195.605 277.305 196.175 ;
  END
 END i230
 PIN i231
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 193.895 277.305 194.465 ;
  END
 END i231
 PIN i232
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 191.235 277.305 191.805 ;
  END
 END i232
 PIN i233
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 189.525 277.305 190.095 ;
  END
 END i233
 PIN i234
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 186.865 277.305 187.435 ;
  END
 END i234
 PIN i235
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 185.155 277.305 185.725 ;
  END
 END i235
 PIN i236
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 182.495 277.305 183.065 ;
  END
 END i236
 PIN i237
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 259.445 277.305 260.015 ;
  END
 END i237
 PIN i238
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 180.785 277.305 181.355 ;
  END
 END i238
 PIN i239
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 178.125 277.305 178.695 ;
  END
 END i239
 PIN i240
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 176.415 277.305 176.985 ;
  END
 END i240
 PIN i241
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 173.755 277.305 174.325 ;
  END
 END i241
 PIN i242
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 172.045 277.305 172.615 ;
  END
 END i242
 PIN i243
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 169.385 277.305 169.955 ;
  END
 END i243
 PIN i244
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 153.615 277.305 154.185 ;
  END
 END i244
 PIN i245
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 150.955 277.305 151.525 ;
  END
 END i245
 PIN i246
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 114.855 277.305 115.425 ;
  END
 END i246
 PIN i247
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 112.195 277.305 112.765 ;
  END
 END i247
 PIN i248
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 256.785 277.305 257.355 ;
  END
 END i248
 PIN i249
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 110.485 277.305 111.055 ;
  END
 END i249
 PIN i250
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 107.825 277.305 108.395 ;
  END
 END i250
 PIN i251
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 106.115 277.305 106.685 ;
  END
 END i251
 PIN i252
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 103.455 277.305 104.025 ;
  END
 END i252
 PIN i253
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 101.745 277.305 102.315 ;
  END
 END i253
 PIN i254
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 99.085 277.305 99.655 ;
  END
 END i254
 PIN i255
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 97.375 277.305 97.945 ;
  END
 END i255
 PIN i256
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 94.715 277.305 95.285 ;
  END
 END i256
 PIN i257
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 93.005 277.305 93.575 ;
  END
 END i257
 PIN i258
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 90.345 277.305 90.915 ;
  END
 END i258
 PIN i259
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 255.075 277.305 255.645 ;
  END
 END i259
 PIN i260
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 88.635 277.305 89.205 ;
  END
 END i260
 PIN i261
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 85.975 277.305 86.545 ;
  END
 END i261
 PIN i262
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 84.265 277.305 84.835 ;
  END
 END i262
 PIN i263
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 81.605 277.305 82.175 ;
  END
 END i263
 PIN i264
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 79.895 277.305 80.465 ;
  END
 END i264
 PIN i265
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 77.235 277.305 77.805 ;
  END
 END i265
 PIN i266
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 75.525 277.305 76.095 ;
  END
 END i266
 PIN i267
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 72.865 277.305 73.435 ;
  END
 END i267
 PIN i268
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 71.155 277.305 71.725 ;
  END
 END i268
 PIN i269
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 68.495 277.305 69.065 ;
  END
 END i269
 PIN i270
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 252.415 277.305 252.985 ;
  END
 END i270
 PIN i271
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 66.785 277.305 67.355 ;
  END
 END i271
 PIN i272
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 64.125 277.305 64.695 ;
  END
 END i272
 PIN i273
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 62.415 277.305 62.985 ;
  END
 END i273
 PIN i274
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 59.755 277.305 60.325 ;
  END
 END i274
 PIN i275
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 58.045 277.305 58.615 ;
  END
 END i275
 PIN i276
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 55.385 277.305 55.955 ;
  END
 END i276
 PIN i277
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 53.675 277.305 54.245 ;
  END
 END i277
 PIN i278
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 51.015 277.305 51.585 ;
  END
 END i278
 PIN i279
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 49.305 277.305 49.875 ;
  END
 END i279
 PIN i280
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 46.645 277.305 47.215 ;
  END
 END i280
 PIN i281
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 250.705 277.305 251.275 ;
  END
 END i281
 PIN i282
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 44.935 277.305 45.505 ;
  END
 END i282
 PIN i283
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 42.275 277.305 42.845 ;
  END
 END i283
 PIN i284
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 40.565 277.305 41.135 ;
  END
 END i284
 PIN i285
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 37.905 277.305 38.475 ;
  END
 END i285
 PIN i286
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 36.195 277.305 36.765 ;
  END
 END i286
 PIN i287
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 33.535 277.305 34.105 ;
  END
 END i287
 PIN i288
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 31.825 277.305 32.395 ;
  END
 END i288
 PIN i289
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 29.165 277.305 29.735 ;
  END
 END i289
 PIN i290
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 27.455 277.305 28.025 ;
  END
 END i290
 PIN i291
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 24.795 277.305 25.365 ;
  END
 END i291
 PIN i292
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 248.045 277.305 248.615 ;
  END
 END i292
 PIN i293
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 23.085 277.305 23.655 ;
  END
 END i293
 PIN i294
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 20.425 277.305 20.995 ;
  END
 END i294
 PIN i295
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 283.575 277.305 284.145 ;
  END
 END i295
 PIN i296
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 134.615 277.305 135.185 ;
  END
 END i296
 PIN i297
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 302.955 276.545 303.525 ;
  END
 END i297
 PIN i298
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 299.345 276.545 299.915 ;
  END
 END i298
 PIN i299
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 246.715 276.545 247.285 ;
  END
 END i299
 PIN i300
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 243.105 276.545 243.675 ;
  END
 END i300
 PIN i301
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 242.345 276.545 242.915 ;
  END
 END i301
 PIN i302
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 238.735 276.545 239.305 ;
  END
 END i302
 PIN i303
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 237.975 276.545 238.545 ;
  END
 END i303
 PIN i304
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 234.365 276.545 234.935 ;
  END
 END i304
 PIN i305
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 233.605 276.545 234.175 ;
  END
 END i305
 PIN i306
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 229.995 276.545 230.565 ;
  END
 END i306
 PIN i307
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 229.235 276.545 229.805 ;
  END
 END i307
 PIN i308
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 225.625 276.545 226.195 ;
  END
 END i308
 PIN i309
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 264.195 276.545 264.765 ;
  END
 END i309
 PIN i310
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 224.865 276.545 225.435 ;
  END
 END i310
 PIN i311
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 221.255 276.545 221.825 ;
  END
 END i311
 PIN i312
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 220.495 276.545 221.065 ;
  END
 END i312
 PIN i313
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 216.885 276.545 217.455 ;
  END
 END i313
 PIN i314
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 216.125 276.545 216.695 ;
  END
 END i314
 PIN i315
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 212.515 276.545 213.085 ;
  END
 END i315
 PIN i316
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 211.755 276.545 212.325 ;
  END
 END i316
 PIN i317
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 208.145 276.545 208.715 ;
  END
 END i317
 PIN i318
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 207.385 276.545 207.955 ;
  END
 END i318
 PIN i319
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 203.775 276.545 204.345 ;
  END
 END i319
 PIN i320
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 260.585 276.545 261.155 ;
  END
 END i320
 PIN i321
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 203.015 276.545 203.585 ;
  END
 END i321
 PIN i322
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 199.405 276.545 199.975 ;
  END
 END i322
 PIN i323
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 198.645 276.545 199.215 ;
  END
 END i323
 PIN i324
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 195.035 276.545 195.605 ;
  END
 END i324
 PIN i325
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 194.275 276.545 194.845 ;
  END
 END i325
 PIN i326
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 190.665 276.545 191.235 ;
  END
 END i326
 PIN i327
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 189.905 276.545 190.475 ;
  END
 END i327
 PIN i328
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 186.295 276.545 186.865 ;
  END
 END i328
 PIN i329
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 185.535 276.545 186.105 ;
  END
 END i329
 PIN i330
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 181.925 276.545 182.495 ;
  END
 END i330
 PIN i331
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 259.825 276.545 260.395 ;
  END
 END i331
 PIN i332
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 181.165 276.545 181.735 ;
  END
 END i332
 PIN i333
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 177.555 276.545 178.125 ;
  END
 END i333
 PIN i334
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 176.795 276.545 177.365 ;
  END
 END i334
 PIN i335
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 173.185 276.545 173.755 ;
  END
 END i335
 PIN i336
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 172.425 276.545 172.995 ;
  END
 END i336
 PIN i337
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 168.815 276.545 169.385 ;
  END
 END i337
 PIN i338
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 154.185 276.545 154.755 ;
  END
 END i338
 PIN i339
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 150.575 276.545 151.145 ;
  END
 END i339
 PIN i340
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 115.235 276.545 115.805 ;
  END
 END i340
 PIN i341
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 111.625 276.545 112.195 ;
  END
 END i341
 PIN i342
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 256.215 276.545 256.785 ;
  END
 END i342
 PIN i343
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 110.865 276.545 111.435 ;
  END
 END i343
 PIN i344
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 107.255 276.545 107.825 ;
  END
 END i344
 PIN i345
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 106.495 276.545 107.065 ;
  END
 END i345
 PIN i346
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 102.885 276.545 103.455 ;
  END
 END i346
 PIN i347
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 102.125 276.545 102.695 ;
  END
 END i347
 PIN i348
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 98.515 276.545 99.085 ;
  END
 END i348
 PIN i349
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 97.755 276.545 98.325 ;
  END
 END i349
 PIN i350
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 94.145 276.545 94.715 ;
  END
 END i350
 PIN i351
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 93.385 276.545 93.955 ;
  END
 END i351
 PIN i352
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 89.775 276.545 90.345 ;
  END
 END i352
 PIN i353
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 255.455 276.545 256.025 ;
  END
 END i353
 PIN i354
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 89.015 276.545 89.585 ;
  END
 END i354
 PIN i355
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 85.405 276.545 85.975 ;
  END
 END i355
 PIN i356
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 84.645 276.545 85.215 ;
  END
 END i356
 PIN i357
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 81.035 276.545 81.605 ;
  END
 END i357
 PIN i358
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 80.275 276.545 80.845 ;
  END
 END i358
 PIN i359
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 76.665 276.545 77.235 ;
  END
 END i359
 PIN i360
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 75.905 276.545 76.475 ;
  END
 END i360
 PIN i361
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 72.295 276.545 72.865 ;
  END
 END i361
 PIN i362
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 71.535 276.545 72.105 ;
  END
 END i362
 PIN i363
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 67.925 276.545 68.495 ;
  END
 END i363
 PIN i364
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 251.845 276.545 252.415 ;
  END
 END i364
 PIN i365
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 67.165 276.545 67.735 ;
  END
 END i365
 PIN i366
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 63.555 276.545 64.125 ;
  END
 END i366
 PIN i367
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 62.795 276.545 63.365 ;
  END
 END i367
 PIN i368
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 59.185 276.545 59.755 ;
  END
 END i368
 PIN i369
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 58.425 276.545 58.995 ;
  END
 END i369
 PIN i370
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 54.815 276.545 55.385 ;
  END
 END i370
 PIN i371
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 54.055 276.545 54.625 ;
  END
 END i371
 PIN i372
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 50.445 276.545 51.015 ;
  END
 END i372
 PIN i373
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 49.685 276.545 50.255 ;
  END
 END i373
 PIN i374
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 46.075 276.545 46.645 ;
  END
 END i374
 PIN i375
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 251.085 276.545 251.655 ;
  END
 END i375
 PIN i376
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 45.315 276.545 45.885 ;
  END
 END i376
 PIN i377
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 41.705 276.545 42.275 ;
  END
 END i377
 PIN i378
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 40.945 276.545 41.515 ;
  END
 END i378
 PIN i379
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 37.335 276.545 37.905 ;
  END
 END i379
 PIN i380
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 36.575 276.545 37.145 ;
  END
 END i380
 PIN i381
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 32.965 276.545 33.535 ;
  END
 END i381
 PIN i382
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 32.205 276.545 32.775 ;
  END
 END i382
 PIN i383
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 28.595 276.545 29.165 ;
  END
 END i383
 PIN i384
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 27.835 276.545 28.405 ;
  END
 END i384
 PIN i385
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 24.225 276.545 24.795 ;
  END
 END i385
 PIN i386
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 247.475 276.545 248.045 ;
  END
 END i386
 PIN i387
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 23.465 276.545 24.035 ;
  END
 END i387
 PIN i388
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 19.855 276.545 20.425 ;
  END
 END i388
 PIN i389
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 210.235 348.365 210.805 348.935 ;
  END
 END i389
 PIN i390
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 215.555 348.365 216.125 348.935 ;
  END
 END i390
 PIN i391
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 214.795 348.365 215.365 348.935 ;
  END
 END i391
 PIN i392
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 214.035 348.365 214.605 348.935 ;
  END
 END i392
 PIN i393
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 212.895 348.365 213.465 348.935 ;
  END
 END i393
 PIN i394
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 212.135 348.365 212.705 348.935 ;
  END
 END i394
 PIN i395
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 210.995 348.365 211.565 348.935 ;
  END
 END i395
 PIN i396
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 204.915 348.365 205.485 348.935 ;
  END
 END i396
 PIN i397
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 234.555 348.365 235.125 348.935 ;
  END
 END i397
 PIN i398
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 225.815 348.365 226.385 348.935 ;
  END
 END i398
 PIN i399
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 233.415 348.365 233.985 348.935 ;
  END
 END i399
 PIN i400
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 226.575 348.365 227.145 348.935 ;
  END
 END i400
 PIN i401
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 232.655 348.365 233.225 348.935 ;
  END
 END i401
 PIN i402
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 227.715 348.365 228.285 348.935 ;
  END
 END i402
 PIN i403
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 178.315 348.365 178.885 348.935 ;
  END
 END i403
 PIN i404
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 348.365 175.465 348.935 ;
  END
 END i404
 PIN i405
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 159.315 348.365 159.885 348.935 ;
  END
 END i405
 PIN i406
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.755 348.365 155.325 348.935 ;
  END
 END i406
 PIN i407
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 152.855 348.365 153.425 348.935 ;
  END
 END i407
 PIN i408
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 150.195 348.365 150.765 348.935 ;
  END
 END i408
 PIN i409
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 148.295 348.365 148.865 348.935 ;
  END
 END i409
 PIN i410
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 183.635 348.365 184.205 348.935 ;
  END
 END i410
 PIN i411
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 186.675 348.365 187.245 348.935 ;
  END
 END i411
 PIN i412
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 189.335 348.365 189.905 348.935 ;
  END
 END i412
 PIN i413
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 193.895 348.365 194.465 348.935 ;
  END
 END i413
 PIN i414
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 160.075 348.365 160.645 348.935 ;
  END
 END i414
 PIN i415
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 170.335 348.365 170.905 348.935 ;
  END
 END i415
 PIN i416
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 166.535 348.365 167.105 348.935 ;
  END
 END i416
 PIN i417
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 162.735 348.365 163.305 348.935 ;
  END
 END i417
 PIN i418
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 167.295 348.365 167.865 348.935 ;
  END
 END i418
 PIN i419
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 171.095 348.365 171.665 348.935 ;
  END
 END i419
 PIN i420
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 348.365 176.225 348.935 ;
  END
 END i420
 PIN i421
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 179.455 348.365 180.025 348.935 ;
  END
 END i421
 PIN i422
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 163.875 348.365 164.445 348.935 ;
  END
 END i422
 PIN i423
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 201.495 348.365 202.065 348.935 ;
  END
 END i423
 PIN i424
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 200.355 348.365 200.925 348.935 ;
  END
 END i424
 PIN i425
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 197.695 348.365 198.265 348.935 ;
  END
 END i425
 PIN i426
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 196.555 348.365 197.125 348.935 ;
  END
 END i426
 PIN i427
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 193.135 348.365 193.705 348.935 ;
  END
 END i427
 PIN i428
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 191.995 348.365 192.565 348.935 ;
  END
 END i428
 PIN i429
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 190.475 348.365 191.045 348.935 ;
  END
 END i429
 PIN i430
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.395 348.365 203.965 348.935 ;
  END
 END i430
 OBS
  LAYER metal1 ;
   RECT 0 0 280.06 350.55 ;
  LAYER via1 ;
   RECT 0 0 280.06 350.55 ;
  LAYER metal2 ;
   RECT 0 0 280.06 350.55 ;
  LAYER via2 ;
   RECT 0 0 280.06 350.55 ;
  LAYER metal3 ;
   RECT 0 0 280.06 350.55 ;
  LAYER via3 ;
   RECT 0 0 280.06 350.55 ;
  LAYER metal4 ;
   RECT 0 0 280.06 350.55 ;
 END
END block_737x1845_682

MACRO block_644x666_92
 CLASS BLOCK ;
 FOREIGN block_644x666_92 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 244.72 BY 126.54 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 33.535 241.585 34.105 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 33.915 240.825 34.485 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 34.295 241.585 34.865 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 34.675 240.825 35.245 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 35.055 241.585 35.625 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 35.435 240.825 36.005 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 35.815 241.585 36.385 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 36.195 240.825 36.765 ;
  END
 END o7
 PIN o8
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 36.575 241.585 37.145 ;
  END
 END o8
 PIN o9
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 36.955 240.825 37.525 ;
  END
 END o9
 PIN o10
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 38.095 241.585 38.665 ;
  END
 END o10
 PIN o11
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 38.475 240.825 39.045 ;
  END
 END o11
 PIN o12
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 38.855 241.585 39.425 ;
  END
 END o12
 PIN o13
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 39.235 240.825 39.805 ;
  END
 END o13
 PIN o14
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 39.615 241.585 40.185 ;
  END
 END o14
 PIN o15
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 39.995 240.825 40.565 ;
  END
 END o15
 PIN o16
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 40.375 241.585 40.945 ;
  END
 END o16
 PIN o17
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 40.755 240.825 41.325 ;
  END
 END o17
 PIN o18
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 41.135 241.585 41.705 ;
  END
 END o18
 PIN o19
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 43.415 241.585 43.985 ;
  END
 END o19
 PIN o20
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 43.795 240.825 44.365 ;
  END
 END o20
 PIN o21
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 44.175 241.585 44.745 ;
  END
 END o21
 PIN o22
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 44.555 240.825 45.125 ;
  END
 END o22
 PIN o23
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 44.935 241.585 45.505 ;
  END
 END o23
 PIN o24
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 45.315 240.825 45.885 ;
  END
 END o24
 PIN o25
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 45.695 241.585 46.265 ;
  END
 END o25
 PIN o26
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 46.075 240.825 46.645 ;
  END
 END o26
 PIN o27
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 47.215 241.585 47.785 ;
  END
 END o27
 PIN o28
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 47.595 240.825 48.165 ;
  END
 END o28
 PIN o29
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 47.975 241.585 48.545 ;
  END
 END o29
 PIN o30
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 177.175 86.45 177.745 87.02 ;
  END
 END o30
 PIN o31
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 49.495 241.585 50.065 ;
  END
 END o31
 PIN o32
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 49.875 240.825 50.445 ;
  END
 END o32
 PIN o33
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 50.255 241.585 50.825 ;
  END
 END o33
 PIN o34
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 68.115 241.585 68.685 ;
  END
 END o34
 PIN o35
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 68.875 241.585 69.445 ;
  END
 END o35
 PIN o36
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 70.395 241.585 70.965 ;
  END
 END o36
 PIN o37
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 70.775 240.825 71.345 ;
  END
 END o37
 PIN o38
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 71.155 241.585 71.725 ;
  END
 END o38
 PIN o39
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 71.535 240.825 72.105 ;
  END
 END o39
 PIN o40
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 50.635 240.825 51.205 ;
  END
 END o40
 PIN o41
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 52.535 241.585 53.105 ;
  END
 END o41
 PIN o42
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 52.915 240.825 53.485 ;
  END
 END o42
 PIN o43
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 53.675 241.585 54.245 ;
  END
 END o43
 PIN o44
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 54.055 240.825 54.625 ;
  END
 END o44
 PIN o45
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 54.435 241.585 55.005 ;
  END
 END o45
 PIN o46
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 54.815 240.825 55.385 ;
  END
 END o46
 PIN o47
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 55.195 241.585 55.765 ;
  END
 END o47
 PIN o48
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 56.335 241.585 56.905 ;
  END
 END o48
 PIN o49
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 56.715 240.825 57.285 ;
  END
 END o49
 PIN o50
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 57.095 241.585 57.665 ;
  END
 END o50
 PIN o51
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 57.475 240.825 58.045 ;
  END
 END o51
 PIN o52
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 57.855 241.585 58.425 ;
  END
 END o52
 PIN o53
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 58.235 240.825 58.805 ;
  END
 END o53
 PIN o54
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 58.615 241.585 59.185 ;
  END
 END o54
 PIN o55
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 58.995 240.825 59.565 ;
  END
 END o55
 PIN o56
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 59.375 241.585 59.945 ;
  END
 END o56
 PIN o57
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 59.755 240.825 60.325 ;
  END
 END o57
 PIN o58
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 63.935 124.545 64.505 125.115 ;
  END
 END o58
 PIN o59
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 67.355 124.545 67.925 125.115 ;
  END
 END o59
 PIN o60
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 80.655 124.545 81.225 125.115 ;
  END
 END o60
 PIN o61
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 98.515 124.545 99.085 125.115 ;
  END
 END o61
 PIN o62
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 48.355 3.325 48.925 ;
  END
 END o62
 PIN o63
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 40.375 3.325 40.945 ;
  END
 END o63
 PIN o64
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 39.615 3.325 40.185 ;
  END
 END o64
 PIN o65
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 47.975 4.085 48.545 ;
  END
 END o65
 PIN o66
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 44.935 3.325 45.505 ;
  END
 END o66
 PIN o67
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 44.175 3.325 44.745 ;
  END
 END o67
 PIN o68
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 124.545 130.245 125.115 ;
  END
 END o68
 PIN o69
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 135.375 124.545 135.945 125.115 ;
  END
 END o69
 PIN o70
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 168.435 124.545 169.005 125.115 ;
  END
 END o70
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 37.335 124.545 37.905 125.115 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 33.915 124.545 34.485 125.115 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 36.195 124.545 36.765 125.115 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 43.795 124.545 44.365 125.115 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 51.775 124.545 52.345 125.115 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 52.915 124.545 53.485 125.115 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 54.815 124.545 55.385 125.115 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 56.335 124.545 56.905 125.115 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 57.475 124.545 58.045 125.115 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 59.375 124.545 59.945 125.115 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 60.515 124.545 61.085 125.115 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 47.215 124.545 47.785 125.115 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 49.495 124.545 50.065 125.115 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 48.355 124.545 48.925 125.115 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 60.895 241.585 61.465 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 65.075 124.545 65.645 125.115 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 63.935 241.585 64.505 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 96.235 124.545 96.805 125.115 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 63.935 3.325 64.505 ;
  END
 END i18
 PIN i19
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 127.395 124.545 127.965 125.115 ;
  END
 END i19
 PIN i20
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 166.155 124.545 166.725 125.115 ;
  END
 END i20
 OBS
  LAYER metal1 ;
   RECT 0 0 244.72 126.54 ;
  LAYER via1 ;
   RECT 0 0 244.72 126.54 ;
  LAYER metal2 ;
   RECT 0 0 244.72 126.54 ;
  LAYER via2 ;
   RECT 0 0 244.72 126.54 ;
  LAYER metal3 ;
   RECT 0 0 244.72 126.54 ;
  LAYER via3 ;
   RECT 0 0 244.72 126.54 ;
  LAYER metal4 ;
   RECT 0 0 244.72 126.54 ;
 END
END block_644x666_92

MACRO block_321x315_66
 CLASS BLOCK ;
 FOREIGN block_321x315_66 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 121.98 BY 59.85 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 48.735 3.325 49.305 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 44.175 118.845 44.745 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 34.295 3.325 34.865 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 35.815 3.325 36.385 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 38.095 3.325 38.665 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 39.615 3.325 40.185 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 41.135 3.325 41.705 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 42.655 3.325 43.225 ;
  END
 END o7
 PIN o8
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 44.175 3.325 44.745 ;
  END
 END o8
 PIN o9
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 45.695 3.325 46.265 ;
  END
 END o9
 PIN o10
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 22.895 118.845 23.465 ;
  END
 END o10
 PIN o11
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 6.935 3.325 7.505 ;
  END
 END o11
 PIN o12
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 7.695 3.325 8.265 ;
  END
 END o12
 PIN o13
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 19.855 3.325 20.425 ;
  END
 END o13
 PIN o14
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 21.375 3.325 21.945 ;
  END
 END o14
 PIN o15
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 22.135 3.325 22.705 ;
  END
 END o15
 PIN o16
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 24.415 3.325 24.985 ;
  END
 END o16
 PIN o17
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 25.935 3.325 26.505 ;
  END
 END o17
 PIN o18
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 26.695 3.325 27.265 ;
  END
 END o18
 PIN o19
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 27.455 3.325 28.025 ;
  END
 END o19
 PIN o20
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 28.975 3.325 29.545 ;
  END
 END o20
 PIN o21
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 30.495 3.325 31.065 ;
  END
 END o21
 PIN o22
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 32.015 3.325 32.585 ;
  END
 END o22
 PIN o23
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 9.215 3.325 9.785 ;
  END
 END o23
 PIN o24
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 10.735 3.325 11.305 ;
  END
 END o24
 PIN o25
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 11.495 3.325 12.065 ;
  END
 END o25
 PIN o26
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 12.255 3.325 12.825 ;
  END
 END o26
 PIN o27
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 13.775 3.325 14.345 ;
  END
 END o27
 PIN o28
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 15.295 3.325 15.865 ;
  END
 END o28
 PIN o29
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 16.055 3.325 16.625 ;
  END
 END o29
 PIN o30
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 16.815 3.325 17.385 ;
  END
 END o30
 PIN o31
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 25.175 118.845 25.745 ;
  END
 END o31
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 32.015 118.845 32.585 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 44.935 118.845 45.505 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 30.495 118.845 31.065 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 31.255 118.845 31.825 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 35.055 118.845 35.625 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 34.295 118.845 34.865 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 27.455 118.845 28.025 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 28.975 118.845 29.545 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 24.415 118.845 24.985 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 42.655 118.845 43.225 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 47.215 3.325 47.785 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 4.655 3.325 5.225 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 22.135 118.845 22.705 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 21.375 118.845 21.945 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 29.735 118.845 30.305 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 26.695 118.845 27.265 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 25.935 118.845 26.505 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 3.895 118.845 4.465 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 4.655 118.845 5.225 ;
  END
 END i18
 PIN i19
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 6.175 118.845 6.745 ;
  END
 END i19
 PIN i20
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 6.935 118.845 7.505 ;
  END
 END i20
 PIN i21
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 7.695 118.845 8.265 ;
  END
 END i21
 PIN i22
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 8.455 118.845 9.025 ;
  END
 END i22
 PIN i23
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 9.215 118.845 9.785 ;
  END
 END i23
 PIN i24
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 10.735 118.845 11.305 ;
  END
 END i24
 PIN i25
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 11.495 118.845 12.065 ;
  END
 END i25
 PIN i26
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 12.255 118.845 12.825 ;
  END
 END i26
 PIN i27
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 13.015 118.845 13.585 ;
  END
 END i27
 PIN i28
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 13.775 118.845 14.345 ;
  END
 END i28
 PIN i29
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 15.295 118.845 15.865 ;
  END
 END i29
 PIN i30
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 16.055 118.845 16.625 ;
  END
 END i30
 PIN i31
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 16.815 118.845 17.385 ;
  END
 END i31
 PIN i32
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 17.575 118.845 18.145 ;
  END
 END i32
 PIN i33
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 18.335 118.845 18.905 ;
  END
 END i33
 OBS
  LAYER metal1 ;
   RECT 0 0 121.98 59.85 ;
  LAYER via1 ;
   RECT 0 0 121.98 59.85 ;
  LAYER metal2 ;
   RECT 0 0 121.98 59.85 ;
  LAYER via2 ;
   RECT 0 0 121.98 59.85 ;
  LAYER metal3 ;
   RECT 0 0 121.98 59.85 ;
  LAYER via3 ;
   RECT 0 0 121.98 59.85 ;
  LAYER metal4 ;
   RECT 0 0 121.98 59.85 ;
 END
END block_321x315_66

MACRO block_779x1431_153
 CLASS BLOCK ;
 FOREIGN block_779x1431_153 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 296.02 BY 271.89 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 4.275 269.325 4.845 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 12.445 269.325 13.015 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 104.215 269.325 104.785 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 112.385 269.325 112.955 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 120.555 269.325 121.125 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 157.035 269.325 157.605 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 165.205 269.325 165.775 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 173.375 269.325 173.945 ;
  END
 END o7
 PIN o8
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 181.545 269.325 182.115 ;
  END
 END o8
 PIN o9
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 189.715 269.325 190.285 ;
  END
 END o9
 PIN o10
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 197.885 269.325 198.455 ;
  END
 END o10
 PIN o11
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 224.295 269.325 224.865 ;
  END
 END o11
 PIN o12
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 20.615 269.325 21.185 ;
  END
 END o12
 PIN o13
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 232.465 269.325 233.035 ;
  END
 END o13
 PIN o14
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 240.635 269.325 241.205 ;
  END
 END o14
 PIN o15
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 248.805 269.325 249.375 ;
  END
 END o15
 PIN o16
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 256.975 269.325 257.545 ;
  END
 END o16
 PIN o17
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 265.145 269.325 265.715 ;
  END
 END o17
 PIN o18
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 28.785 269.325 29.355 ;
  END
 END o18
 PIN o19
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 36.955 269.325 37.525 ;
  END
 END o19
 PIN o20
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 45.125 269.325 45.695 ;
  END
 END o20
 PIN o21
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 53.295 269.325 53.865 ;
  END
 END o21
 PIN o22
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 79.705 269.325 80.275 ;
  END
 END o22
 PIN o23
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 87.875 269.325 88.445 ;
  END
 END o23
 PIN o24
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 96.045 269.325 96.615 ;
  END
 END o24
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 291.935 127.585 292.505 128.155 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 291.935 144.685 292.505 145.255 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 291.935 132.905 292.505 133.475 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 291.935 137.275 292.505 137.845 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 291.175 127.965 291.745 128.535 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 291.175 127.205 291.745 127.775 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 291.935 126.825 292.505 127.395 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 291.935 136.515 292.505 137.085 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 291.935 149.625 292.505 150.195 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 291.175 144.305 291.745 144.875 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 291.935 141.075 292.505 141.645 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 291.935 143.925 292.505 144.495 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 291.935 146.015 292.505 146.585 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 291.935 148.485 292.505 149.055 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 291.175 150.005 291.745 150.575 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 282.435 126.445 283.005 127.015 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 282.435 139.745 283.005 140.315 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 2.565 269.325 3.135 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 10.735 269.325 11.305 ;
  END
 END i18
 PIN i19
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 102.505 269.325 103.075 ;
  END
 END i19
 PIN i20
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 110.675 269.325 111.245 ;
  END
 END i20
 PIN i21
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 118.845 269.325 119.415 ;
  END
 END i21
 PIN i22
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 158.745 269.325 159.315 ;
  END
 END i22
 PIN i23
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 166.915 269.325 167.485 ;
  END
 END i23
 PIN i24
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 175.085 269.325 175.655 ;
  END
 END i24
 PIN i25
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 183.255 269.325 183.825 ;
  END
 END i25
 PIN i26
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 191.425 269.325 191.995 ;
  END
 END i26
 PIN i27
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 199.595 269.325 200.165 ;
  END
 END i27
 PIN i28
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 226.005 269.325 226.575 ;
  END
 END i28
 PIN i29
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 18.905 269.325 19.475 ;
  END
 END i29
 PIN i30
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 234.175 269.325 234.745 ;
  END
 END i30
 PIN i31
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 242.345 269.325 242.915 ;
  END
 END i31
 PIN i32
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 250.515 269.325 251.085 ;
  END
 END i32
 PIN i33
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 258.685 269.325 259.255 ;
  END
 END i33
 PIN i34
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 266.855 269.325 267.425 ;
  END
 END i34
 PIN i35
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 27.075 269.325 27.645 ;
  END
 END i35
 PIN i36
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 35.245 269.325 35.815 ;
  END
 END i36
 PIN i37
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 43.415 269.325 43.985 ;
  END
 END i37
 PIN i38
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 51.585 269.325 52.155 ;
  END
 END i38
 PIN i39
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 77.995 269.325 78.565 ;
  END
 END i39
 PIN i40
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 86.165 269.325 86.735 ;
  END
 END i40
 PIN i41
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 94.335 269.325 94.905 ;
  END
 END i41
 PIN i42
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 33.535 269.325 34.105 ;
  END
 END i42
 PIN i43
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 37.525 268.565 38.095 ;
  END
 END i43
 PIN i44
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 41.705 269.325 42.275 ;
  END
 END i44
 PIN i45
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 25.365 269.325 25.935 ;
  END
 END i45
 PIN i46
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 100.795 269.325 101.365 ;
  END
 END i46
 PIN i47
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 104.785 268.565 105.355 ;
  END
 END i47
 PIN i48
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 108.965 269.325 109.535 ;
  END
 END i48
 PIN i49
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 112.955 268.565 113.525 ;
  END
 END i49
 PIN i50
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 176.795 269.325 177.365 ;
  END
 END i50
 PIN i51
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 172.805 268.565 173.375 ;
  END
 END i51
 PIN i52
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 168.625 269.325 169.195 ;
  END
 END i52
 PIN i53
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 164.635 268.565 165.205 ;
  END
 END i53
 PIN i54
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 244.055 269.325 244.625 ;
  END
 END i54
 PIN i55
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 240.065 268.565 240.635 ;
  END
 END i55
 PIN i56
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 235.885 269.325 236.455 ;
  END
 END i56
 PIN i57
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 252.225 269.325 252.795 ;
  END
 END i57
 PIN i58
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 29.355 268.565 29.925 ;
  END
 END i58
 PIN i59
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 96.615 268.565 97.185 ;
  END
 END i59
 PIN i60
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 180.975 268.565 181.545 ;
  END
 END i60
 PIN i61
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 248.235 268.565 248.805 ;
  END
 END i61
 PIN i62
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 277.115 126.445 277.685 127.015 ;
  END
 END i62
 PIN i63
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 277.115 139.745 277.685 140.315 ;
  END
 END i63
 PIN i64
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 3.135 268.565 3.705 ;
  END
 END i64
 PIN i65
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 11.305 268.565 11.875 ;
  END
 END i65
 PIN i66
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 103.075 268.565 103.645 ;
  END
 END i66
 PIN i67
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 111.245 268.565 111.815 ;
  END
 END i67
 PIN i68
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 119.415 268.565 119.985 ;
  END
 END i68
 PIN i69
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 158.175 268.565 158.745 ;
  END
 END i69
 PIN i70
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 166.345 268.565 166.915 ;
  END
 END i70
 PIN i71
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 174.515 268.565 175.085 ;
  END
 END i71
 PIN i72
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 182.685 268.565 183.255 ;
  END
 END i72
 PIN i73
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 190.855 268.565 191.425 ;
  END
 END i73
 PIN i74
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 199.025 268.565 199.595 ;
  END
 END i74
 PIN i75
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 225.435 268.565 226.005 ;
  END
 END i75
 PIN i76
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 19.475 268.565 20.045 ;
  END
 END i76
 PIN i77
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 233.605 268.565 234.175 ;
  END
 END i77
 PIN i78
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 241.775 268.565 242.345 ;
  END
 END i78
 PIN i79
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 249.945 268.565 250.515 ;
  END
 END i79
 PIN i80
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 258.115 268.565 258.685 ;
  END
 END i80
 PIN i81
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 266.285 268.565 266.855 ;
  END
 END i81
 PIN i82
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 27.645 268.565 28.215 ;
  END
 END i82
 PIN i83
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 35.815 268.565 36.385 ;
  END
 END i83
 PIN i84
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 43.985 268.565 44.555 ;
  END
 END i84
 PIN i85
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 52.155 268.565 52.725 ;
  END
 END i85
 PIN i86
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 78.565 268.565 79.135 ;
  END
 END i86
 PIN i87
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 86.735 268.565 87.305 ;
  END
 END i87
 PIN i88
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 94.905 268.565 95.475 ;
  END
 END i88
 PIN i89
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 291.935 134.045 292.505 134.615 ;
  END
 END i89
 PIN i90
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 291.175 134.425 291.745 134.995 ;
  END
 END i90
 PIN i91
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.235 3.705 267.805 4.275 ;
  END
 END i91
 PIN i92
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.235 11.875 267.805 12.445 ;
  END
 END i92
 PIN i93
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.235 103.645 267.805 104.215 ;
  END
 END i93
 PIN i94
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.235 111.815 267.805 112.385 ;
  END
 END i94
 PIN i95
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.235 119.985 267.805 120.555 ;
  END
 END i95
 PIN i96
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.235 157.605 267.805 158.175 ;
  END
 END i96
 PIN i97
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.235 165.775 267.805 166.345 ;
  END
 END i97
 PIN i98
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.235 173.945 267.805 174.515 ;
  END
 END i98
 PIN i99
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.235 182.115 267.805 182.685 ;
  END
 END i99
 PIN i100
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.235 190.285 267.805 190.855 ;
  END
 END i100
 PIN i101
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.235 198.455 267.805 199.025 ;
  END
 END i101
 PIN i102
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.235 224.865 267.805 225.435 ;
  END
 END i102
 PIN i103
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.235 20.045 267.805 20.615 ;
  END
 END i103
 PIN i104
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.235 233.035 267.805 233.605 ;
  END
 END i104
 PIN i105
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.235 241.205 267.805 241.775 ;
  END
 END i105
 PIN i106
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.235 249.375 267.805 249.945 ;
  END
 END i106
 PIN i107
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.235 257.545 267.805 258.115 ;
  END
 END i107
 PIN i108
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.235 265.715 267.805 266.285 ;
  END
 END i108
 PIN i109
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.235 28.215 267.805 28.785 ;
  END
 END i109
 PIN i110
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.235 36.385 267.805 36.955 ;
  END
 END i110
 PIN i111
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.235 44.555 267.805 45.125 ;
  END
 END i111
 PIN i112
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.235 52.725 267.805 53.295 ;
  END
 END i112
 PIN i113
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.235 79.135 267.805 79.705 ;
  END
 END i113
 PIN i114
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.235 87.305 267.805 87.875 ;
  END
 END i114
 PIN i115
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.235 95.475 267.805 96.045 ;
  END
 END i115
 PIN i116
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 291.175 126.445 291.745 127.015 ;
  END
 END i116
 PIN i117
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 290.035 126.445 290.605 127.015 ;
  END
 END i117
 PIN i118
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 288.135 126.445 288.705 127.015 ;
  END
 END i118
 PIN i119
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 286.615 126.445 287.185 127.015 ;
  END
 END i119
 PIN i120
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 285.095 126.445 285.665 127.015 ;
  END
 END i120
 PIN i121
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 283.195 126.445 283.765 127.015 ;
  END
 END i121
 PIN i122
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 291.175 139.745 291.745 140.315 ;
  END
 END i122
 PIN i123
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 290.035 139.745 290.605 140.315 ;
  END
 END i123
 PIN i124
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 288.135 139.745 288.705 140.315 ;
  END
 END i124
 PIN i125
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 286.615 139.745 287.185 140.315 ;
  END
 END i125
 PIN i126
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 285.095 139.745 285.665 140.315 ;
  END
 END i126
 PIN i127
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 283.195 139.745 283.765 140.315 ;
  END
 END i127
 OBS
  LAYER metal1 ;
   RECT 0.0 0.0 272.84 1.71 ;
   RECT 0.0 1.71 272.84 3.42 ;
   RECT 0.0 3.42 272.84 5.13 ;
   RECT 0.0 5.13 272.84 6.84 ;
   RECT 0.0 6.84 272.84 8.55 ;
   RECT 0.0 8.55 272.84 10.26 ;
   RECT 0.0 10.26 272.84 11.97 ;
   RECT 0.0 11.97 272.84 13.68 ;
   RECT 0.0 13.68 272.84 15.39 ;
   RECT 0.0 15.39 272.84 17.1 ;
   RECT 0.0 17.1 272.84 18.81 ;
   RECT 0.0 18.81 272.84 20.52 ;
   RECT 0.0 20.52 272.84 22.23 ;
   RECT 0.0 22.23 272.84 23.94 ;
   RECT 0.0 23.94 272.84 25.65 ;
   RECT 0.0 25.65 272.84 27.36 ;
   RECT 0.0 27.36 272.84 29.07 ;
   RECT 0.0 29.07 272.84 30.78 ;
   RECT 0.0 30.78 272.84 32.49 ;
   RECT 0.0 32.49 272.84 34.2 ;
   RECT 0.0 34.2 272.84 35.91 ;
   RECT 0.0 35.91 272.84 37.62 ;
   RECT 0.0 37.62 272.84 39.33 ;
   RECT 0.0 39.33 272.84 41.04 ;
   RECT 0.0 41.04 272.84 42.75 ;
   RECT 0.0 42.75 272.84 44.46 ;
   RECT 0.0 44.46 272.84 46.17 ;
   RECT 0.0 46.17 272.84 47.88 ;
   RECT 0.0 47.88 272.84 49.59 ;
   RECT 0.0 49.59 272.84 51.3 ;
   RECT 0.0 51.3 272.84 53.01 ;
   RECT 0.0 53.01 272.84 54.72 ;
   RECT 0.0 54.72 272.84 56.43 ;
   RECT 0.0 56.43 272.84 58.14 ;
   RECT 0.0 58.14 272.84 59.85 ;
   RECT 0.0 59.85 272.84 61.56 ;
   RECT 0.0 61.56 272.84 63.27 ;
   RECT 0.0 63.27 272.84 64.98 ;
   RECT 0.0 64.98 272.84 66.69 ;
   RECT 0.0 66.69 272.84 68.4 ;
   RECT 0.0 68.4 272.84 70.11 ;
   RECT 0.0 70.11 272.84 71.82 ;
   RECT 0.0 71.82 272.84 73.53 ;
   RECT 0.0 73.53 272.84 75.24 ;
   RECT 0.0 75.24 272.84 76.95 ;
   RECT 0.0 76.95 272.84 78.66 ;
   RECT 0.0 78.66 272.84 80.37 ;
   RECT 0.0 80.37 272.84 82.08 ;
   RECT 0.0 82.08 272.84 83.79 ;
   RECT 0.0 83.79 272.84 85.5 ;
   RECT 0.0 85.5 272.84 87.21 ;
   RECT 0.0 87.21 272.84 88.92 ;
   RECT 0.0 88.92 272.84 90.63 ;
   RECT 0.0 90.63 272.84 92.34 ;
   RECT 0.0 92.34 272.84 94.05 ;
   RECT 0.0 94.05 272.84 95.76 ;
   RECT 0.0 95.76 272.84 97.47 ;
   RECT 0.0 97.47 272.84 99.18 ;
   RECT 0.0 99.18 272.84 100.89 ;
   RECT 0.0 100.89 272.84 102.6 ;
   RECT 0.0 102.6 272.84 104.31 ;
   RECT 0.0 104.31 272.84 106.02 ;
   RECT 0.0 106.02 272.84 107.73 ;
   RECT 0.0 107.73 272.84 109.44 ;
   RECT 0.0 109.44 272.84 111.15 ;
   RECT 0.0 111.15 272.84 112.86 ;
   RECT 0.0 112.86 272.84 114.57 ;
   RECT 0.0 114.57 272.84 116.28 ;
   RECT 0.0 116.28 272.84 117.99 ;
   RECT 0.0 117.99 272.84 119.7 ;
   RECT 0.0 119.7 272.84 121.41 ;
   RECT 0.0 121.41 272.84 123.12 ;
   RECT 0.0 123.12 272.84 124.83 ;
   RECT 0.0 124.83 296.02 126.54 ;
   RECT 0.0 126.54 296.02 128.25 ;
   RECT 0.0 128.25 296.02 129.96 ;
   RECT 0.0 129.96 296.02 131.67 ;
   RECT 0.0 131.67 296.02 133.38 ;
   RECT 0.0 133.38 296.02 135.09 ;
   RECT 0.0 135.09 296.02 136.8 ;
   RECT 0.0 136.8 296.02 138.51 ;
   RECT 0.0 138.51 296.02 140.22 ;
   RECT 0.0 140.22 296.02 141.93 ;
   RECT 0.0 141.93 296.02 143.64 ;
   RECT 0.0 143.64 296.02 145.35 ;
   RECT 0.0 145.35 296.02 147.06 ;
   RECT 0.0 147.06 296.02 148.77 ;
   RECT 0.0 148.77 296.02 150.48 ;
   RECT 0.0 150.48 296.02 152.19 ;
   RECT 0.0 152.19 296.02 153.9 ;
   RECT 0.0 153.9 272.84 155.61 ;
   RECT 0.0 155.61 272.84 157.32 ;
   RECT 0.0 157.32 272.84 159.03 ;
   RECT 0.0 159.03 272.84 160.74 ;
   RECT 0.0 160.74 272.84 162.45 ;
   RECT 0.0 162.45 272.84 164.16 ;
   RECT 0.0 164.16 272.84 165.87 ;
   RECT 0.0 165.87 272.84 167.58 ;
   RECT 0.0 167.58 272.84 169.29 ;
   RECT 0.0 169.29 272.84 171.0 ;
   RECT 0.0 171.0 272.84 172.71 ;
   RECT 0.0 172.71 272.84 174.42 ;
   RECT 0.0 174.42 272.84 176.13 ;
   RECT 0.0 176.13 272.84 177.84 ;
   RECT 0.0 177.84 272.84 179.55 ;
   RECT 0.0 179.55 272.84 181.26 ;
   RECT 0.0 181.26 272.84 182.97 ;
   RECT 0.0 182.97 272.84 184.68 ;
   RECT 0.0 184.68 272.84 186.39 ;
   RECT 0.0 186.39 272.84 188.1 ;
   RECT 0.0 188.1 272.84 189.81 ;
   RECT 0.0 189.81 272.84 191.52 ;
   RECT 0.0 191.52 272.84 193.23 ;
   RECT 0.0 193.23 272.84 194.94 ;
   RECT 0.0 194.94 272.84 196.65 ;
   RECT 0.0 196.65 272.84 198.36 ;
   RECT 0.0 198.36 272.84 200.07 ;
   RECT 0.0 200.07 272.84 201.78 ;
   RECT 0.0 201.78 272.84 203.49 ;
   RECT 0.0 203.49 272.84 205.2 ;
   RECT 0.0 205.2 272.84 206.91 ;
   RECT 0.0 206.91 272.84 208.62 ;
   RECT 0.0 208.62 272.84 210.33 ;
   RECT 0.0 210.33 272.84 212.04 ;
   RECT 0.0 212.04 272.84 213.75 ;
   RECT 0.0 213.75 272.84 215.46 ;
   RECT 0.0 215.46 272.84 217.17 ;
   RECT 0.0 217.17 272.84 218.88 ;
   RECT 0.0 218.88 272.84 220.59 ;
   RECT 0.0 220.59 272.84 222.3 ;
   RECT 0.0 222.3 272.84 224.01 ;
   RECT 0.0 224.01 272.84 225.72 ;
   RECT 0.0 225.72 272.84 227.43 ;
   RECT 0.0 227.43 272.84 229.14 ;
   RECT 0.0 229.14 272.84 230.85 ;
   RECT 0.0 230.85 272.84 232.56 ;
   RECT 0.0 232.56 272.84 234.27 ;
   RECT 0.0 234.27 272.84 235.98 ;
   RECT 0.0 235.98 272.84 237.69 ;
   RECT 0.0 237.69 272.84 239.4 ;
   RECT 0.0 239.4 272.84 241.11 ;
   RECT 0.0 241.11 272.84 242.82 ;
   RECT 0.0 242.82 272.84 244.53 ;
   RECT 0.0 244.53 272.84 246.24 ;
   RECT 0.0 246.24 272.84 247.95 ;
   RECT 0.0 247.95 272.84 249.66 ;
   RECT 0.0 249.66 272.84 251.37 ;
   RECT 0.0 251.37 272.84 253.08 ;
   RECT 0.0 253.08 272.84 254.79 ;
   RECT 0.0 254.79 272.84 256.5 ;
   RECT 0.0 256.5 272.84 258.21 ;
   RECT 0.0 258.21 272.84 259.92 ;
   RECT 0.0 259.92 272.84 261.63 ;
   RECT 0.0 261.63 272.84 263.34 ;
   RECT 0.0 263.34 272.84 265.05 ;
   RECT 0.0 265.05 272.84 266.76 ;
   RECT 0.0 266.76 272.84 268.47 ;
   RECT 0.0 268.47 272.84 270.18 ;
   RECT 0.0 270.18 272.84 271.89 ;
  LAYER via1 ;
   RECT 0.0 0.0 272.84 1.71 ;
   RECT 0.0 1.71 272.84 3.42 ;
   RECT 0.0 3.42 272.84 5.13 ;
   RECT 0.0 5.13 272.84 6.84 ;
   RECT 0.0 6.84 272.84 8.55 ;
   RECT 0.0 8.55 272.84 10.26 ;
   RECT 0.0 10.26 272.84 11.97 ;
   RECT 0.0 11.97 272.84 13.68 ;
   RECT 0.0 13.68 272.84 15.39 ;
   RECT 0.0 15.39 272.84 17.1 ;
   RECT 0.0 17.1 272.84 18.81 ;
   RECT 0.0 18.81 272.84 20.52 ;
   RECT 0.0 20.52 272.84 22.23 ;
   RECT 0.0 22.23 272.84 23.94 ;
   RECT 0.0 23.94 272.84 25.65 ;
   RECT 0.0 25.65 272.84 27.36 ;
   RECT 0.0 27.36 272.84 29.07 ;
   RECT 0.0 29.07 272.84 30.78 ;
   RECT 0.0 30.78 272.84 32.49 ;
   RECT 0.0 32.49 272.84 34.2 ;
   RECT 0.0 34.2 272.84 35.91 ;
   RECT 0.0 35.91 272.84 37.62 ;
   RECT 0.0 37.62 272.84 39.33 ;
   RECT 0.0 39.33 272.84 41.04 ;
   RECT 0.0 41.04 272.84 42.75 ;
   RECT 0.0 42.75 272.84 44.46 ;
   RECT 0.0 44.46 272.84 46.17 ;
   RECT 0.0 46.17 272.84 47.88 ;
   RECT 0.0 47.88 272.84 49.59 ;
   RECT 0.0 49.59 272.84 51.3 ;
   RECT 0.0 51.3 272.84 53.01 ;
   RECT 0.0 53.01 272.84 54.72 ;
   RECT 0.0 54.72 272.84 56.43 ;
   RECT 0.0 56.43 272.84 58.14 ;
   RECT 0.0 58.14 272.84 59.85 ;
   RECT 0.0 59.85 272.84 61.56 ;
   RECT 0.0 61.56 272.84 63.27 ;
   RECT 0.0 63.27 272.84 64.98 ;
   RECT 0.0 64.98 272.84 66.69 ;
   RECT 0.0 66.69 272.84 68.4 ;
   RECT 0.0 68.4 272.84 70.11 ;
   RECT 0.0 70.11 272.84 71.82 ;
   RECT 0.0 71.82 272.84 73.53 ;
   RECT 0.0 73.53 272.84 75.24 ;
   RECT 0.0 75.24 272.84 76.95 ;
   RECT 0.0 76.95 272.84 78.66 ;
   RECT 0.0 78.66 272.84 80.37 ;
   RECT 0.0 80.37 272.84 82.08 ;
   RECT 0.0 82.08 272.84 83.79 ;
   RECT 0.0 83.79 272.84 85.5 ;
   RECT 0.0 85.5 272.84 87.21 ;
   RECT 0.0 87.21 272.84 88.92 ;
   RECT 0.0 88.92 272.84 90.63 ;
   RECT 0.0 90.63 272.84 92.34 ;
   RECT 0.0 92.34 272.84 94.05 ;
   RECT 0.0 94.05 272.84 95.76 ;
   RECT 0.0 95.76 272.84 97.47 ;
   RECT 0.0 97.47 272.84 99.18 ;
   RECT 0.0 99.18 272.84 100.89 ;
   RECT 0.0 100.89 272.84 102.6 ;
   RECT 0.0 102.6 272.84 104.31 ;
   RECT 0.0 104.31 272.84 106.02 ;
   RECT 0.0 106.02 272.84 107.73 ;
   RECT 0.0 107.73 272.84 109.44 ;
   RECT 0.0 109.44 272.84 111.15 ;
   RECT 0.0 111.15 272.84 112.86 ;
   RECT 0.0 112.86 272.84 114.57 ;
   RECT 0.0 114.57 272.84 116.28 ;
   RECT 0.0 116.28 272.84 117.99 ;
   RECT 0.0 117.99 272.84 119.7 ;
   RECT 0.0 119.7 272.84 121.41 ;
   RECT 0.0 121.41 272.84 123.12 ;
   RECT 0.0 123.12 272.84 124.83 ;
   RECT 0.0 124.83 296.02 126.54 ;
   RECT 0.0 126.54 296.02 128.25 ;
   RECT 0.0 128.25 296.02 129.96 ;
   RECT 0.0 129.96 296.02 131.67 ;
   RECT 0.0 131.67 296.02 133.38 ;
   RECT 0.0 133.38 296.02 135.09 ;
   RECT 0.0 135.09 296.02 136.8 ;
   RECT 0.0 136.8 296.02 138.51 ;
   RECT 0.0 138.51 296.02 140.22 ;
   RECT 0.0 140.22 296.02 141.93 ;
   RECT 0.0 141.93 296.02 143.64 ;
   RECT 0.0 143.64 296.02 145.35 ;
   RECT 0.0 145.35 296.02 147.06 ;
   RECT 0.0 147.06 296.02 148.77 ;
   RECT 0.0 148.77 296.02 150.48 ;
   RECT 0.0 150.48 296.02 152.19 ;
   RECT 0.0 152.19 296.02 153.9 ;
   RECT 0.0 153.9 272.84 155.61 ;
   RECT 0.0 155.61 272.84 157.32 ;
   RECT 0.0 157.32 272.84 159.03 ;
   RECT 0.0 159.03 272.84 160.74 ;
   RECT 0.0 160.74 272.84 162.45 ;
   RECT 0.0 162.45 272.84 164.16 ;
   RECT 0.0 164.16 272.84 165.87 ;
   RECT 0.0 165.87 272.84 167.58 ;
   RECT 0.0 167.58 272.84 169.29 ;
   RECT 0.0 169.29 272.84 171.0 ;
   RECT 0.0 171.0 272.84 172.71 ;
   RECT 0.0 172.71 272.84 174.42 ;
   RECT 0.0 174.42 272.84 176.13 ;
   RECT 0.0 176.13 272.84 177.84 ;
   RECT 0.0 177.84 272.84 179.55 ;
   RECT 0.0 179.55 272.84 181.26 ;
   RECT 0.0 181.26 272.84 182.97 ;
   RECT 0.0 182.97 272.84 184.68 ;
   RECT 0.0 184.68 272.84 186.39 ;
   RECT 0.0 186.39 272.84 188.1 ;
   RECT 0.0 188.1 272.84 189.81 ;
   RECT 0.0 189.81 272.84 191.52 ;
   RECT 0.0 191.52 272.84 193.23 ;
   RECT 0.0 193.23 272.84 194.94 ;
   RECT 0.0 194.94 272.84 196.65 ;
   RECT 0.0 196.65 272.84 198.36 ;
   RECT 0.0 198.36 272.84 200.07 ;
   RECT 0.0 200.07 272.84 201.78 ;
   RECT 0.0 201.78 272.84 203.49 ;
   RECT 0.0 203.49 272.84 205.2 ;
   RECT 0.0 205.2 272.84 206.91 ;
   RECT 0.0 206.91 272.84 208.62 ;
   RECT 0.0 208.62 272.84 210.33 ;
   RECT 0.0 210.33 272.84 212.04 ;
   RECT 0.0 212.04 272.84 213.75 ;
   RECT 0.0 213.75 272.84 215.46 ;
   RECT 0.0 215.46 272.84 217.17 ;
   RECT 0.0 217.17 272.84 218.88 ;
   RECT 0.0 218.88 272.84 220.59 ;
   RECT 0.0 220.59 272.84 222.3 ;
   RECT 0.0 222.3 272.84 224.01 ;
   RECT 0.0 224.01 272.84 225.72 ;
   RECT 0.0 225.72 272.84 227.43 ;
   RECT 0.0 227.43 272.84 229.14 ;
   RECT 0.0 229.14 272.84 230.85 ;
   RECT 0.0 230.85 272.84 232.56 ;
   RECT 0.0 232.56 272.84 234.27 ;
   RECT 0.0 234.27 272.84 235.98 ;
   RECT 0.0 235.98 272.84 237.69 ;
   RECT 0.0 237.69 272.84 239.4 ;
   RECT 0.0 239.4 272.84 241.11 ;
   RECT 0.0 241.11 272.84 242.82 ;
   RECT 0.0 242.82 272.84 244.53 ;
   RECT 0.0 244.53 272.84 246.24 ;
   RECT 0.0 246.24 272.84 247.95 ;
   RECT 0.0 247.95 272.84 249.66 ;
   RECT 0.0 249.66 272.84 251.37 ;
   RECT 0.0 251.37 272.84 253.08 ;
   RECT 0.0 253.08 272.84 254.79 ;
   RECT 0.0 254.79 272.84 256.5 ;
   RECT 0.0 256.5 272.84 258.21 ;
   RECT 0.0 258.21 272.84 259.92 ;
   RECT 0.0 259.92 272.84 261.63 ;
   RECT 0.0 261.63 272.84 263.34 ;
   RECT 0.0 263.34 272.84 265.05 ;
   RECT 0.0 265.05 272.84 266.76 ;
   RECT 0.0 266.76 272.84 268.47 ;
   RECT 0.0 268.47 272.84 270.18 ;
   RECT 0.0 270.18 272.84 271.89 ;
  LAYER metal2 ;
   RECT 0.0 0.0 272.84 1.71 ;
   RECT 0.0 1.71 272.84 3.42 ;
   RECT 0.0 3.42 272.84 5.13 ;
   RECT 0.0 5.13 272.84 6.84 ;
   RECT 0.0 6.84 272.84 8.55 ;
   RECT 0.0 8.55 272.84 10.26 ;
   RECT 0.0 10.26 272.84 11.97 ;
   RECT 0.0 11.97 272.84 13.68 ;
   RECT 0.0 13.68 272.84 15.39 ;
   RECT 0.0 15.39 272.84 17.1 ;
   RECT 0.0 17.1 272.84 18.81 ;
   RECT 0.0 18.81 272.84 20.52 ;
   RECT 0.0 20.52 272.84 22.23 ;
   RECT 0.0 22.23 272.84 23.94 ;
   RECT 0.0 23.94 272.84 25.65 ;
   RECT 0.0 25.65 272.84 27.36 ;
   RECT 0.0 27.36 272.84 29.07 ;
   RECT 0.0 29.07 272.84 30.78 ;
   RECT 0.0 30.78 272.84 32.49 ;
   RECT 0.0 32.49 272.84 34.2 ;
   RECT 0.0 34.2 272.84 35.91 ;
   RECT 0.0 35.91 272.84 37.62 ;
   RECT 0.0 37.62 272.84 39.33 ;
   RECT 0.0 39.33 272.84 41.04 ;
   RECT 0.0 41.04 272.84 42.75 ;
   RECT 0.0 42.75 272.84 44.46 ;
   RECT 0.0 44.46 272.84 46.17 ;
   RECT 0.0 46.17 272.84 47.88 ;
   RECT 0.0 47.88 272.84 49.59 ;
   RECT 0.0 49.59 272.84 51.3 ;
   RECT 0.0 51.3 272.84 53.01 ;
   RECT 0.0 53.01 272.84 54.72 ;
   RECT 0.0 54.72 272.84 56.43 ;
   RECT 0.0 56.43 272.84 58.14 ;
   RECT 0.0 58.14 272.84 59.85 ;
   RECT 0.0 59.85 272.84 61.56 ;
   RECT 0.0 61.56 272.84 63.27 ;
   RECT 0.0 63.27 272.84 64.98 ;
   RECT 0.0 64.98 272.84 66.69 ;
   RECT 0.0 66.69 272.84 68.4 ;
   RECT 0.0 68.4 272.84 70.11 ;
   RECT 0.0 70.11 272.84 71.82 ;
   RECT 0.0 71.82 272.84 73.53 ;
   RECT 0.0 73.53 272.84 75.24 ;
   RECT 0.0 75.24 272.84 76.95 ;
   RECT 0.0 76.95 272.84 78.66 ;
   RECT 0.0 78.66 272.84 80.37 ;
   RECT 0.0 80.37 272.84 82.08 ;
   RECT 0.0 82.08 272.84 83.79 ;
   RECT 0.0 83.79 272.84 85.5 ;
   RECT 0.0 85.5 272.84 87.21 ;
   RECT 0.0 87.21 272.84 88.92 ;
   RECT 0.0 88.92 272.84 90.63 ;
   RECT 0.0 90.63 272.84 92.34 ;
   RECT 0.0 92.34 272.84 94.05 ;
   RECT 0.0 94.05 272.84 95.76 ;
   RECT 0.0 95.76 272.84 97.47 ;
   RECT 0.0 97.47 272.84 99.18 ;
   RECT 0.0 99.18 272.84 100.89 ;
   RECT 0.0 100.89 272.84 102.6 ;
   RECT 0.0 102.6 272.84 104.31 ;
   RECT 0.0 104.31 272.84 106.02 ;
   RECT 0.0 106.02 272.84 107.73 ;
   RECT 0.0 107.73 272.84 109.44 ;
   RECT 0.0 109.44 272.84 111.15 ;
   RECT 0.0 111.15 272.84 112.86 ;
   RECT 0.0 112.86 272.84 114.57 ;
   RECT 0.0 114.57 272.84 116.28 ;
   RECT 0.0 116.28 272.84 117.99 ;
   RECT 0.0 117.99 272.84 119.7 ;
   RECT 0.0 119.7 272.84 121.41 ;
   RECT 0.0 121.41 272.84 123.12 ;
   RECT 0.0 123.12 272.84 124.83 ;
   RECT 0.0 124.83 296.02 126.54 ;
   RECT 0.0 126.54 296.02 128.25 ;
   RECT 0.0 128.25 296.02 129.96 ;
   RECT 0.0 129.96 296.02 131.67 ;
   RECT 0.0 131.67 296.02 133.38 ;
   RECT 0.0 133.38 296.02 135.09 ;
   RECT 0.0 135.09 296.02 136.8 ;
   RECT 0.0 136.8 296.02 138.51 ;
   RECT 0.0 138.51 296.02 140.22 ;
   RECT 0.0 140.22 296.02 141.93 ;
   RECT 0.0 141.93 296.02 143.64 ;
   RECT 0.0 143.64 296.02 145.35 ;
   RECT 0.0 145.35 296.02 147.06 ;
   RECT 0.0 147.06 296.02 148.77 ;
   RECT 0.0 148.77 296.02 150.48 ;
   RECT 0.0 150.48 296.02 152.19 ;
   RECT 0.0 152.19 296.02 153.9 ;
   RECT 0.0 153.9 272.84 155.61 ;
   RECT 0.0 155.61 272.84 157.32 ;
   RECT 0.0 157.32 272.84 159.03 ;
   RECT 0.0 159.03 272.84 160.74 ;
   RECT 0.0 160.74 272.84 162.45 ;
   RECT 0.0 162.45 272.84 164.16 ;
   RECT 0.0 164.16 272.84 165.87 ;
   RECT 0.0 165.87 272.84 167.58 ;
   RECT 0.0 167.58 272.84 169.29 ;
   RECT 0.0 169.29 272.84 171.0 ;
   RECT 0.0 171.0 272.84 172.71 ;
   RECT 0.0 172.71 272.84 174.42 ;
   RECT 0.0 174.42 272.84 176.13 ;
   RECT 0.0 176.13 272.84 177.84 ;
   RECT 0.0 177.84 272.84 179.55 ;
   RECT 0.0 179.55 272.84 181.26 ;
   RECT 0.0 181.26 272.84 182.97 ;
   RECT 0.0 182.97 272.84 184.68 ;
   RECT 0.0 184.68 272.84 186.39 ;
   RECT 0.0 186.39 272.84 188.1 ;
   RECT 0.0 188.1 272.84 189.81 ;
   RECT 0.0 189.81 272.84 191.52 ;
   RECT 0.0 191.52 272.84 193.23 ;
   RECT 0.0 193.23 272.84 194.94 ;
   RECT 0.0 194.94 272.84 196.65 ;
   RECT 0.0 196.65 272.84 198.36 ;
   RECT 0.0 198.36 272.84 200.07 ;
   RECT 0.0 200.07 272.84 201.78 ;
   RECT 0.0 201.78 272.84 203.49 ;
   RECT 0.0 203.49 272.84 205.2 ;
   RECT 0.0 205.2 272.84 206.91 ;
   RECT 0.0 206.91 272.84 208.62 ;
   RECT 0.0 208.62 272.84 210.33 ;
   RECT 0.0 210.33 272.84 212.04 ;
   RECT 0.0 212.04 272.84 213.75 ;
   RECT 0.0 213.75 272.84 215.46 ;
   RECT 0.0 215.46 272.84 217.17 ;
   RECT 0.0 217.17 272.84 218.88 ;
   RECT 0.0 218.88 272.84 220.59 ;
   RECT 0.0 220.59 272.84 222.3 ;
   RECT 0.0 222.3 272.84 224.01 ;
   RECT 0.0 224.01 272.84 225.72 ;
   RECT 0.0 225.72 272.84 227.43 ;
   RECT 0.0 227.43 272.84 229.14 ;
   RECT 0.0 229.14 272.84 230.85 ;
   RECT 0.0 230.85 272.84 232.56 ;
   RECT 0.0 232.56 272.84 234.27 ;
   RECT 0.0 234.27 272.84 235.98 ;
   RECT 0.0 235.98 272.84 237.69 ;
   RECT 0.0 237.69 272.84 239.4 ;
   RECT 0.0 239.4 272.84 241.11 ;
   RECT 0.0 241.11 272.84 242.82 ;
   RECT 0.0 242.82 272.84 244.53 ;
   RECT 0.0 244.53 272.84 246.24 ;
   RECT 0.0 246.24 272.84 247.95 ;
   RECT 0.0 247.95 272.84 249.66 ;
   RECT 0.0 249.66 272.84 251.37 ;
   RECT 0.0 251.37 272.84 253.08 ;
   RECT 0.0 253.08 272.84 254.79 ;
   RECT 0.0 254.79 272.84 256.5 ;
   RECT 0.0 256.5 272.84 258.21 ;
   RECT 0.0 258.21 272.84 259.92 ;
   RECT 0.0 259.92 272.84 261.63 ;
   RECT 0.0 261.63 272.84 263.34 ;
   RECT 0.0 263.34 272.84 265.05 ;
   RECT 0.0 265.05 272.84 266.76 ;
   RECT 0.0 266.76 272.84 268.47 ;
   RECT 0.0 268.47 272.84 270.18 ;
   RECT 0.0 270.18 272.84 271.89 ;
  LAYER via2 ;
   RECT 0.0 0.0 272.84 1.71 ;
   RECT 0.0 1.71 272.84 3.42 ;
   RECT 0.0 3.42 272.84 5.13 ;
   RECT 0.0 5.13 272.84 6.84 ;
   RECT 0.0 6.84 272.84 8.55 ;
   RECT 0.0 8.55 272.84 10.26 ;
   RECT 0.0 10.26 272.84 11.97 ;
   RECT 0.0 11.97 272.84 13.68 ;
   RECT 0.0 13.68 272.84 15.39 ;
   RECT 0.0 15.39 272.84 17.1 ;
   RECT 0.0 17.1 272.84 18.81 ;
   RECT 0.0 18.81 272.84 20.52 ;
   RECT 0.0 20.52 272.84 22.23 ;
   RECT 0.0 22.23 272.84 23.94 ;
   RECT 0.0 23.94 272.84 25.65 ;
   RECT 0.0 25.65 272.84 27.36 ;
   RECT 0.0 27.36 272.84 29.07 ;
   RECT 0.0 29.07 272.84 30.78 ;
   RECT 0.0 30.78 272.84 32.49 ;
   RECT 0.0 32.49 272.84 34.2 ;
   RECT 0.0 34.2 272.84 35.91 ;
   RECT 0.0 35.91 272.84 37.62 ;
   RECT 0.0 37.62 272.84 39.33 ;
   RECT 0.0 39.33 272.84 41.04 ;
   RECT 0.0 41.04 272.84 42.75 ;
   RECT 0.0 42.75 272.84 44.46 ;
   RECT 0.0 44.46 272.84 46.17 ;
   RECT 0.0 46.17 272.84 47.88 ;
   RECT 0.0 47.88 272.84 49.59 ;
   RECT 0.0 49.59 272.84 51.3 ;
   RECT 0.0 51.3 272.84 53.01 ;
   RECT 0.0 53.01 272.84 54.72 ;
   RECT 0.0 54.72 272.84 56.43 ;
   RECT 0.0 56.43 272.84 58.14 ;
   RECT 0.0 58.14 272.84 59.85 ;
   RECT 0.0 59.85 272.84 61.56 ;
   RECT 0.0 61.56 272.84 63.27 ;
   RECT 0.0 63.27 272.84 64.98 ;
   RECT 0.0 64.98 272.84 66.69 ;
   RECT 0.0 66.69 272.84 68.4 ;
   RECT 0.0 68.4 272.84 70.11 ;
   RECT 0.0 70.11 272.84 71.82 ;
   RECT 0.0 71.82 272.84 73.53 ;
   RECT 0.0 73.53 272.84 75.24 ;
   RECT 0.0 75.24 272.84 76.95 ;
   RECT 0.0 76.95 272.84 78.66 ;
   RECT 0.0 78.66 272.84 80.37 ;
   RECT 0.0 80.37 272.84 82.08 ;
   RECT 0.0 82.08 272.84 83.79 ;
   RECT 0.0 83.79 272.84 85.5 ;
   RECT 0.0 85.5 272.84 87.21 ;
   RECT 0.0 87.21 272.84 88.92 ;
   RECT 0.0 88.92 272.84 90.63 ;
   RECT 0.0 90.63 272.84 92.34 ;
   RECT 0.0 92.34 272.84 94.05 ;
   RECT 0.0 94.05 272.84 95.76 ;
   RECT 0.0 95.76 272.84 97.47 ;
   RECT 0.0 97.47 272.84 99.18 ;
   RECT 0.0 99.18 272.84 100.89 ;
   RECT 0.0 100.89 272.84 102.6 ;
   RECT 0.0 102.6 272.84 104.31 ;
   RECT 0.0 104.31 272.84 106.02 ;
   RECT 0.0 106.02 272.84 107.73 ;
   RECT 0.0 107.73 272.84 109.44 ;
   RECT 0.0 109.44 272.84 111.15 ;
   RECT 0.0 111.15 272.84 112.86 ;
   RECT 0.0 112.86 272.84 114.57 ;
   RECT 0.0 114.57 272.84 116.28 ;
   RECT 0.0 116.28 272.84 117.99 ;
   RECT 0.0 117.99 272.84 119.7 ;
   RECT 0.0 119.7 272.84 121.41 ;
   RECT 0.0 121.41 272.84 123.12 ;
   RECT 0.0 123.12 272.84 124.83 ;
   RECT 0.0 124.83 296.02 126.54 ;
   RECT 0.0 126.54 296.02 128.25 ;
   RECT 0.0 128.25 296.02 129.96 ;
   RECT 0.0 129.96 296.02 131.67 ;
   RECT 0.0 131.67 296.02 133.38 ;
   RECT 0.0 133.38 296.02 135.09 ;
   RECT 0.0 135.09 296.02 136.8 ;
   RECT 0.0 136.8 296.02 138.51 ;
   RECT 0.0 138.51 296.02 140.22 ;
   RECT 0.0 140.22 296.02 141.93 ;
   RECT 0.0 141.93 296.02 143.64 ;
   RECT 0.0 143.64 296.02 145.35 ;
   RECT 0.0 145.35 296.02 147.06 ;
   RECT 0.0 147.06 296.02 148.77 ;
   RECT 0.0 148.77 296.02 150.48 ;
   RECT 0.0 150.48 296.02 152.19 ;
   RECT 0.0 152.19 296.02 153.9 ;
   RECT 0.0 153.9 272.84 155.61 ;
   RECT 0.0 155.61 272.84 157.32 ;
   RECT 0.0 157.32 272.84 159.03 ;
   RECT 0.0 159.03 272.84 160.74 ;
   RECT 0.0 160.74 272.84 162.45 ;
   RECT 0.0 162.45 272.84 164.16 ;
   RECT 0.0 164.16 272.84 165.87 ;
   RECT 0.0 165.87 272.84 167.58 ;
   RECT 0.0 167.58 272.84 169.29 ;
   RECT 0.0 169.29 272.84 171.0 ;
   RECT 0.0 171.0 272.84 172.71 ;
   RECT 0.0 172.71 272.84 174.42 ;
   RECT 0.0 174.42 272.84 176.13 ;
   RECT 0.0 176.13 272.84 177.84 ;
   RECT 0.0 177.84 272.84 179.55 ;
   RECT 0.0 179.55 272.84 181.26 ;
   RECT 0.0 181.26 272.84 182.97 ;
   RECT 0.0 182.97 272.84 184.68 ;
   RECT 0.0 184.68 272.84 186.39 ;
   RECT 0.0 186.39 272.84 188.1 ;
   RECT 0.0 188.1 272.84 189.81 ;
   RECT 0.0 189.81 272.84 191.52 ;
   RECT 0.0 191.52 272.84 193.23 ;
   RECT 0.0 193.23 272.84 194.94 ;
   RECT 0.0 194.94 272.84 196.65 ;
   RECT 0.0 196.65 272.84 198.36 ;
   RECT 0.0 198.36 272.84 200.07 ;
   RECT 0.0 200.07 272.84 201.78 ;
   RECT 0.0 201.78 272.84 203.49 ;
   RECT 0.0 203.49 272.84 205.2 ;
   RECT 0.0 205.2 272.84 206.91 ;
   RECT 0.0 206.91 272.84 208.62 ;
   RECT 0.0 208.62 272.84 210.33 ;
   RECT 0.0 210.33 272.84 212.04 ;
   RECT 0.0 212.04 272.84 213.75 ;
   RECT 0.0 213.75 272.84 215.46 ;
   RECT 0.0 215.46 272.84 217.17 ;
   RECT 0.0 217.17 272.84 218.88 ;
   RECT 0.0 218.88 272.84 220.59 ;
   RECT 0.0 220.59 272.84 222.3 ;
   RECT 0.0 222.3 272.84 224.01 ;
   RECT 0.0 224.01 272.84 225.72 ;
   RECT 0.0 225.72 272.84 227.43 ;
   RECT 0.0 227.43 272.84 229.14 ;
   RECT 0.0 229.14 272.84 230.85 ;
   RECT 0.0 230.85 272.84 232.56 ;
   RECT 0.0 232.56 272.84 234.27 ;
   RECT 0.0 234.27 272.84 235.98 ;
   RECT 0.0 235.98 272.84 237.69 ;
   RECT 0.0 237.69 272.84 239.4 ;
   RECT 0.0 239.4 272.84 241.11 ;
   RECT 0.0 241.11 272.84 242.82 ;
   RECT 0.0 242.82 272.84 244.53 ;
   RECT 0.0 244.53 272.84 246.24 ;
   RECT 0.0 246.24 272.84 247.95 ;
   RECT 0.0 247.95 272.84 249.66 ;
   RECT 0.0 249.66 272.84 251.37 ;
   RECT 0.0 251.37 272.84 253.08 ;
   RECT 0.0 253.08 272.84 254.79 ;
   RECT 0.0 254.79 272.84 256.5 ;
   RECT 0.0 256.5 272.84 258.21 ;
   RECT 0.0 258.21 272.84 259.92 ;
   RECT 0.0 259.92 272.84 261.63 ;
   RECT 0.0 261.63 272.84 263.34 ;
   RECT 0.0 263.34 272.84 265.05 ;
   RECT 0.0 265.05 272.84 266.76 ;
   RECT 0.0 266.76 272.84 268.47 ;
   RECT 0.0 268.47 272.84 270.18 ;
   RECT 0.0 270.18 272.84 271.89 ;
  LAYER metal3 ;
   RECT 0.0 0.0 272.84 1.71 ;
   RECT 0.0 1.71 272.84 3.42 ;
   RECT 0.0 3.42 272.84 5.13 ;
   RECT 0.0 5.13 272.84 6.84 ;
   RECT 0.0 6.84 272.84 8.55 ;
   RECT 0.0 8.55 272.84 10.26 ;
   RECT 0.0 10.26 272.84 11.97 ;
   RECT 0.0 11.97 272.84 13.68 ;
   RECT 0.0 13.68 272.84 15.39 ;
   RECT 0.0 15.39 272.84 17.1 ;
   RECT 0.0 17.1 272.84 18.81 ;
   RECT 0.0 18.81 272.84 20.52 ;
   RECT 0.0 20.52 272.84 22.23 ;
   RECT 0.0 22.23 272.84 23.94 ;
   RECT 0.0 23.94 272.84 25.65 ;
   RECT 0.0 25.65 272.84 27.36 ;
   RECT 0.0 27.36 272.84 29.07 ;
   RECT 0.0 29.07 272.84 30.78 ;
   RECT 0.0 30.78 272.84 32.49 ;
   RECT 0.0 32.49 272.84 34.2 ;
   RECT 0.0 34.2 272.84 35.91 ;
   RECT 0.0 35.91 272.84 37.62 ;
   RECT 0.0 37.62 272.84 39.33 ;
   RECT 0.0 39.33 272.84 41.04 ;
   RECT 0.0 41.04 272.84 42.75 ;
   RECT 0.0 42.75 272.84 44.46 ;
   RECT 0.0 44.46 272.84 46.17 ;
   RECT 0.0 46.17 272.84 47.88 ;
   RECT 0.0 47.88 272.84 49.59 ;
   RECT 0.0 49.59 272.84 51.3 ;
   RECT 0.0 51.3 272.84 53.01 ;
   RECT 0.0 53.01 272.84 54.72 ;
   RECT 0.0 54.72 272.84 56.43 ;
   RECT 0.0 56.43 272.84 58.14 ;
   RECT 0.0 58.14 272.84 59.85 ;
   RECT 0.0 59.85 272.84 61.56 ;
   RECT 0.0 61.56 272.84 63.27 ;
   RECT 0.0 63.27 272.84 64.98 ;
   RECT 0.0 64.98 272.84 66.69 ;
   RECT 0.0 66.69 272.84 68.4 ;
   RECT 0.0 68.4 272.84 70.11 ;
   RECT 0.0 70.11 272.84 71.82 ;
   RECT 0.0 71.82 272.84 73.53 ;
   RECT 0.0 73.53 272.84 75.24 ;
   RECT 0.0 75.24 272.84 76.95 ;
   RECT 0.0 76.95 272.84 78.66 ;
   RECT 0.0 78.66 272.84 80.37 ;
   RECT 0.0 80.37 272.84 82.08 ;
   RECT 0.0 82.08 272.84 83.79 ;
   RECT 0.0 83.79 272.84 85.5 ;
   RECT 0.0 85.5 272.84 87.21 ;
   RECT 0.0 87.21 272.84 88.92 ;
   RECT 0.0 88.92 272.84 90.63 ;
   RECT 0.0 90.63 272.84 92.34 ;
   RECT 0.0 92.34 272.84 94.05 ;
   RECT 0.0 94.05 272.84 95.76 ;
   RECT 0.0 95.76 272.84 97.47 ;
   RECT 0.0 97.47 272.84 99.18 ;
   RECT 0.0 99.18 272.84 100.89 ;
   RECT 0.0 100.89 272.84 102.6 ;
   RECT 0.0 102.6 272.84 104.31 ;
   RECT 0.0 104.31 272.84 106.02 ;
   RECT 0.0 106.02 272.84 107.73 ;
   RECT 0.0 107.73 272.84 109.44 ;
   RECT 0.0 109.44 272.84 111.15 ;
   RECT 0.0 111.15 272.84 112.86 ;
   RECT 0.0 112.86 272.84 114.57 ;
   RECT 0.0 114.57 272.84 116.28 ;
   RECT 0.0 116.28 272.84 117.99 ;
   RECT 0.0 117.99 272.84 119.7 ;
   RECT 0.0 119.7 272.84 121.41 ;
   RECT 0.0 121.41 272.84 123.12 ;
   RECT 0.0 123.12 272.84 124.83 ;
   RECT 0.0 124.83 296.02 126.54 ;
   RECT 0.0 126.54 296.02 128.25 ;
   RECT 0.0 128.25 296.02 129.96 ;
   RECT 0.0 129.96 296.02 131.67 ;
   RECT 0.0 131.67 296.02 133.38 ;
   RECT 0.0 133.38 296.02 135.09 ;
   RECT 0.0 135.09 296.02 136.8 ;
   RECT 0.0 136.8 296.02 138.51 ;
   RECT 0.0 138.51 296.02 140.22 ;
   RECT 0.0 140.22 296.02 141.93 ;
   RECT 0.0 141.93 296.02 143.64 ;
   RECT 0.0 143.64 296.02 145.35 ;
   RECT 0.0 145.35 296.02 147.06 ;
   RECT 0.0 147.06 296.02 148.77 ;
   RECT 0.0 148.77 296.02 150.48 ;
   RECT 0.0 150.48 296.02 152.19 ;
   RECT 0.0 152.19 296.02 153.9 ;
   RECT 0.0 153.9 272.84 155.61 ;
   RECT 0.0 155.61 272.84 157.32 ;
   RECT 0.0 157.32 272.84 159.03 ;
   RECT 0.0 159.03 272.84 160.74 ;
   RECT 0.0 160.74 272.84 162.45 ;
   RECT 0.0 162.45 272.84 164.16 ;
   RECT 0.0 164.16 272.84 165.87 ;
   RECT 0.0 165.87 272.84 167.58 ;
   RECT 0.0 167.58 272.84 169.29 ;
   RECT 0.0 169.29 272.84 171.0 ;
   RECT 0.0 171.0 272.84 172.71 ;
   RECT 0.0 172.71 272.84 174.42 ;
   RECT 0.0 174.42 272.84 176.13 ;
   RECT 0.0 176.13 272.84 177.84 ;
   RECT 0.0 177.84 272.84 179.55 ;
   RECT 0.0 179.55 272.84 181.26 ;
   RECT 0.0 181.26 272.84 182.97 ;
   RECT 0.0 182.97 272.84 184.68 ;
   RECT 0.0 184.68 272.84 186.39 ;
   RECT 0.0 186.39 272.84 188.1 ;
   RECT 0.0 188.1 272.84 189.81 ;
   RECT 0.0 189.81 272.84 191.52 ;
   RECT 0.0 191.52 272.84 193.23 ;
   RECT 0.0 193.23 272.84 194.94 ;
   RECT 0.0 194.94 272.84 196.65 ;
   RECT 0.0 196.65 272.84 198.36 ;
   RECT 0.0 198.36 272.84 200.07 ;
   RECT 0.0 200.07 272.84 201.78 ;
   RECT 0.0 201.78 272.84 203.49 ;
   RECT 0.0 203.49 272.84 205.2 ;
   RECT 0.0 205.2 272.84 206.91 ;
   RECT 0.0 206.91 272.84 208.62 ;
   RECT 0.0 208.62 272.84 210.33 ;
   RECT 0.0 210.33 272.84 212.04 ;
   RECT 0.0 212.04 272.84 213.75 ;
   RECT 0.0 213.75 272.84 215.46 ;
   RECT 0.0 215.46 272.84 217.17 ;
   RECT 0.0 217.17 272.84 218.88 ;
   RECT 0.0 218.88 272.84 220.59 ;
   RECT 0.0 220.59 272.84 222.3 ;
   RECT 0.0 222.3 272.84 224.01 ;
   RECT 0.0 224.01 272.84 225.72 ;
   RECT 0.0 225.72 272.84 227.43 ;
   RECT 0.0 227.43 272.84 229.14 ;
   RECT 0.0 229.14 272.84 230.85 ;
   RECT 0.0 230.85 272.84 232.56 ;
   RECT 0.0 232.56 272.84 234.27 ;
   RECT 0.0 234.27 272.84 235.98 ;
   RECT 0.0 235.98 272.84 237.69 ;
   RECT 0.0 237.69 272.84 239.4 ;
   RECT 0.0 239.4 272.84 241.11 ;
   RECT 0.0 241.11 272.84 242.82 ;
   RECT 0.0 242.82 272.84 244.53 ;
   RECT 0.0 244.53 272.84 246.24 ;
   RECT 0.0 246.24 272.84 247.95 ;
   RECT 0.0 247.95 272.84 249.66 ;
   RECT 0.0 249.66 272.84 251.37 ;
   RECT 0.0 251.37 272.84 253.08 ;
   RECT 0.0 253.08 272.84 254.79 ;
   RECT 0.0 254.79 272.84 256.5 ;
   RECT 0.0 256.5 272.84 258.21 ;
   RECT 0.0 258.21 272.84 259.92 ;
   RECT 0.0 259.92 272.84 261.63 ;
   RECT 0.0 261.63 272.84 263.34 ;
   RECT 0.0 263.34 272.84 265.05 ;
   RECT 0.0 265.05 272.84 266.76 ;
   RECT 0.0 266.76 272.84 268.47 ;
   RECT 0.0 268.47 272.84 270.18 ;
   RECT 0.0 270.18 272.84 271.89 ;
  LAYER via3 ;
   RECT 0.0 0.0 272.84 1.71 ;
   RECT 0.0 1.71 272.84 3.42 ;
   RECT 0.0 3.42 272.84 5.13 ;
   RECT 0.0 5.13 272.84 6.84 ;
   RECT 0.0 6.84 272.84 8.55 ;
   RECT 0.0 8.55 272.84 10.26 ;
   RECT 0.0 10.26 272.84 11.97 ;
   RECT 0.0 11.97 272.84 13.68 ;
   RECT 0.0 13.68 272.84 15.39 ;
   RECT 0.0 15.39 272.84 17.1 ;
   RECT 0.0 17.1 272.84 18.81 ;
   RECT 0.0 18.81 272.84 20.52 ;
   RECT 0.0 20.52 272.84 22.23 ;
   RECT 0.0 22.23 272.84 23.94 ;
   RECT 0.0 23.94 272.84 25.65 ;
   RECT 0.0 25.65 272.84 27.36 ;
   RECT 0.0 27.36 272.84 29.07 ;
   RECT 0.0 29.07 272.84 30.78 ;
   RECT 0.0 30.78 272.84 32.49 ;
   RECT 0.0 32.49 272.84 34.2 ;
   RECT 0.0 34.2 272.84 35.91 ;
   RECT 0.0 35.91 272.84 37.62 ;
   RECT 0.0 37.62 272.84 39.33 ;
   RECT 0.0 39.33 272.84 41.04 ;
   RECT 0.0 41.04 272.84 42.75 ;
   RECT 0.0 42.75 272.84 44.46 ;
   RECT 0.0 44.46 272.84 46.17 ;
   RECT 0.0 46.17 272.84 47.88 ;
   RECT 0.0 47.88 272.84 49.59 ;
   RECT 0.0 49.59 272.84 51.3 ;
   RECT 0.0 51.3 272.84 53.01 ;
   RECT 0.0 53.01 272.84 54.72 ;
   RECT 0.0 54.72 272.84 56.43 ;
   RECT 0.0 56.43 272.84 58.14 ;
   RECT 0.0 58.14 272.84 59.85 ;
   RECT 0.0 59.85 272.84 61.56 ;
   RECT 0.0 61.56 272.84 63.27 ;
   RECT 0.0 63.27 272.84 64.98 ;
   RECT 0.0 64.98 272.84 66.69 ;
   RECT 0.0 66.69 272.84 68.4 ;
   RECT 0.0 68.4 272.84 70.11 ;
   RECT 0.0 70.11 272.84 71.82 ;
   RECT 0.0 71.82 272.84 73.53 ;
   RECT 0.0 73.53 272.84 75.24 ;
   RECT 0.0 75.24 272.84 76.95 ;
   RECT 0.0 76.95 272.84 78.66 ;
   RECT 0.0 78.66 272.84 80.37 ;
   RECT 0.0 80.37 272.84 82.08 ;
   RECT 0.0 82.08 272.84 83.79 ;
   RECT 0.0 83.79 272.84 85.5 ;
   RECT 0.0 85.5 272.84 87.21 ;
   RECT 0.0 87.21 272.84 88.92 ;
   RECT 0.0 88.92 272.84 90.63 ;
   RECT 0.0 90.63 272.84 92.34 ;
   RECT 0.0 92.34 272.84 94.05 ;
   RECT 0.0 94.05 272.84 95.76 ;
   RECT 0.0 95.76 272.84 97.47 ;
   RECT 0.0 97.47 272.84 99.18 ;
   RECT 0.0 99.18 272.84 100.89 ;
   RECT 0.0 100.89 272.84 102.6 ;
   RECT 0.0 102.6 272.84 104.31 ;
   RECT 0.0 104.31 272.84 106.02 ;
   RECT 0.0 106.02 272.84 107.73 ;
   RECT 0.0 107.73 272.84 109.44 ;
   RECT 0.0 109.44 272.84 111.15 ;
   RECT 0.0 111.15 272.84 112.86 ;
   RECT 0.0 112.86 272.84 114.57 ;
   RECT 0.0 114.57 272.84 116.28 ;
   RECT 0.0 116.28 272.84 117.99 ;
   RECT 0.0 117.99 272.84 119.7 ;
   RECT 0.0 119.7 272.84 121.41 ;
   RECT 0.0 121.41 272.84 123.12 ;
   RECT 0.0 123.12 272.84 124.83 ;
   RECT 0.0 124.83 296.02 126.54 ;
   RECT 0.0 126.54 296.02 128.25 ;
   RECT 0.0 128.25 296.02 129.96 ;
   RECT 0.0 129.96 296.02 131.67 ;
   RECT 0.0 131.67 296.02 133.38 ;
   RECT 0.0 133.38 296.02 135.09 ;
   RECT 0.0 135.09 296.02 136.8 ;
   RECT 0.0 136.8 296.02 138.51 ;
   RECT 0.0 138.51 296.02 140.22 ;
   RECT 0.0 140.22 296.02 141.93 ;
   RECT 0.0 141.93 296.02 143.64 ;
   RECT 0.0 143.64 296.02 145.35 ;
   RECT 0.0 145.35 296.02 147.06 ;
   RECT 0.0 147.06 296.02 148.77 ;
   RECT 0.0 148.77 296.02 150.48 ;
   RECT 0.0 150.48 296.02 152.19 ;
   RECT 0.0 152.19 296.02 153.9 ;
   RECT 0.0 153.9 272.84 155.61 ;
   RECT 0.0 155.61 272.84 157.32 ;
   RECT 0.0 157.32 272.84 159.03 ;
   RECT 0.0 159.03 272.84 160.74 ;
   RECT 0.0 160.74 272.84 162.45 ;
   RECT 0.0 162.45 272.84 164.16 ;
   RECT 0.0 164.16 272.84 165.87 ;
   RECT 0.0 165.87 272.84 167.58 ;
   RECT 0.0 167.58 272.84 169.29 ;
   RECT 0.0 169.29 272.84 171.0 ;
   RECT 0.0 171.0 272.84 172.71 ;
   RECT 0.0 172.71 272.84 174.42 ;
   RECT 0.0 174.42 272.84 176.13 ;
   RECT 0.0 176.13 272.84 177.84 ;
   RECT 0.0 177.84 272.84 179.55 ;
   RECT 0.0 179.55 272.84 181.26 ;
   RECT 0.0 181.26 272.84 182.97 ;
   RECT 0.0 182.97 272.84 184.68 ;
   RECT 0.0 184.68 272.84 186.39 ;
   RECT 0.0 186.39 272.84 188.1 ;
   RECT 0.0 188.1 272.84 189.81 ;
   RECT 0.0 189.81 272.84 191.52 ;
   RECT 0.0 191.52 272.84 193.23 ;
   RECT 0.0 193.23 272.84 194.94 ;
   RECT 0.0 194.94 272.84 196.65 ;
   RECT 0.0 196.65 272.84 198.36 ;
   RECT 0.0 198.36 272.84 200.07 ;
   RECT 0.0 200.07 272.84 201.78 ;
   RECT 0.0 201.78 272.84 203.49 ;
   RECT 0.0 203.49 272.84 205.2 ;
   RECT 0.0 205.2 272.84 206.91 ;
   RECT 0.0 206.91 272.84 208.62 ;
   RECT 0.0 208.62 272.84 210.33 ;
   RECT 0.0 210.33 272.84 212.04 ;
   RECT 0.0 212.04 272.84 213.75 ;
   RECT 0.0 213.75 272.84 215.46 ;
   RECT 0.0 215.46 272.84 217.17 ;
   RECT 0.0 217.17 272.84 218.88 ;
   RECT 0.0 218.88 272.84 220.59 ;
   RECT 0.0 220.59 272.84 222.3 ;
   RECT 0.0 222.3 272.84 224.01 ;
   RECT 0.0 224.01 272.84 225.72 ;
   RECT 0.0 225.72 272.84 227.43 ;
   RECT 0.0 227.43 272.84 229.14 ;
   RECT 0.0 229.14 272.84 230.85 ;
   RECT 0.0 230.85 272.84 232.56 ;
   RECT 0.0 232.56 272.84 234.27 ;
   RECT 0.0 234.27 272.84 235.98 ;
   RECT 0.0 235.98 272.84 237.69 ;
   RECT 0.0 237.69 272.84 239.4 ;
   RECT 0.0 239.4 272.84 241.11 ;
   RECT 0.0 241.11 272.84 242.82 ;
   RECT 0.0 242.82 272.84 244.53 ;
   RECT 0.0 244.53 272.84 246.24 ;
   RECT 0.0 246.24 272.84 247.95 ;
   RECT 0.0 247.95 272.84 249.66 ;
   RECT 0.0 249.66 272.84 251.37 ;
   RECT 0.0 251.37 272.84 253.08 ;
   RECT 0.0 253.08 272.84 254.79 ;
   RECT 0.0 254.79 272.84 256.5 ;
   RECT 0.0 256.5 272.84 258.21 ;
   RECT 0.0 258.21 272.84 259.92 ;
   RECT 0.0 259.92 272.84 261.63 ;
   RECT 0.0 261.63 272.84 263.34 ;
   RECT 0.0 263.34 272.84 265.05 ;
   RECT 0.0 265.05 272.84 266.76 ;
   RECT 0.0 266.76 272.84 268.47 ;
   RECT 0.0 268.47 272.84 270.18 ;
   RECT 0.0 270.18 272.84 271.89 ;
  LAYER metal4 ;
   RECT 0.0 0.0 272.84 1.71 ;
   RECT 0.0 1.71 272.84 3.42 ;
   RECT 0.0 3.42 272.84 5.13 ;
   RECT 0.0 5.13 272.84 6.84 ;
   RECT 0.0 6.84 272.84 8.55 ;
   RECT 0.0 8.55 272.84 10.26 ;
   RECT 0.0 10.26 272.84 11.97 ;
   RECT 0.0 11.97 272.84 13.68 ;
   RECT 0.0 13.68 272.84 15.39 ;
   RECT 0.0 15.39 272.84 17.1 ;
   RECT 0.0 17.1 272.84 18.81 ;
   RECT 0.0 18.81 272.84 20.52 ;
   RECT 0.0 20.52 272.84 22.23 ;
   RECT 0.0 22.23 272.84 23.94 ;
   RECT 0.0 23.94 272.84 25.65 ;
   RECT 0.0 25.65 272.84 27.36 ;
   RECT 0.0 27.36 272.84 29.07 ;
   RECT 0.0 29.07 272.84 30.78 ;
   RECT 0.0 30.78 272.84 32.49 ;
   RECT 0.0 32.49 272.84 34.2 ;
   RECT 0.0 34.2 272.84 35.91 ;
   RECT 0.0 35.91 272.84 37.62 ;
   RECT 0.0 37.62 272.84 39.33 ;
   RECT 0.0 39.33 272.84 41.04 ;
   RECT 0.0 41.04 272.84 42.75 ;
   RECT 0.0 42.75 272.84 44.46 ;
   RECT 0.0 44.46 272.84 46.17 ;
   RECT 0.0 46.17 272.84 47.88 ;
   RECT 0.0 47.88 272.84 49.59 ;
   RECT 0.0 49.59 272.84 51.3 ;
   RECT 0.0 51.3 272.84 53.01 ;
   RECT 0.0 53.01 272.84 54.72 ;
   RECT 0.0 54.72 272.84 56.43 ;
   RECT 0.0 56.43 272.84 58.14 ;
   RECT 0.0 58.14 272.84 59.85 ;
   RECT 0.0 59.85 272.84 61.56 ;
   RECT 0.0 61.56 272.84 63.27 ;
   RECT 0.0 63.27 272.84 64.98 ;
   RECT 0.0 64.98 272.84 66.69 ;
   RECT 0.0 66.69 272.84 68.4 ;
   RECT 0.0 68.4 272.84 70.11 ;
   RECT 0.0 70.11 272.84 71.82 ;
   RECT 0.0 71.82 272.84 73.53 ;
   RECT 0.0 73.53 272.84 75.24 ;
   RECT 0.0 75.24 272.84 76.95 ;
   RECT 0.0 76.95 272.84 78.66 ;
   RECT 0.0 78.66 272.84 80.37 ;
   RECT 0.0 80.37 272.84 82.08 ;
   RECT 0.0 82.08 272.84 83.79 ;
   RECT 0.0 83.79 272.84 85.5 ;
   RECT 0.0 85.5 272.84 87.21 ;
   RECT 0.0 87.21 272.84 88.92 ;
   RECT 0.0 88.92 272.84 90.63 ;
   RECT 0.0 90.63 272.84 92.34 ;
   RECT 0.0 92.34 272.84 94.05 ;
   RECT 0.0 94.05 272.84 95.76 ;
   RECT 0.0 95.76 272.84 97.47 ;
   RECT 0.0 97.47 272.84 99.18 ;
   RECT 0.0 99.18 272.84 100.89 ;
   RECT 0.0 100.89 272.84 102.6 ;
   RECT 0.0 102.6 272.84 104.31 ;
   RECT 0.0 104.31 272.84 106.02 ;
   RECT 0.0 106.02 272.84 107.73 ;
   RECT 0.0 107.73 272.84 109.44 ;
   RECT 0.0 109.44 272.84 111.15 ;
   RECT 0.0 111.15 272.84 112.86 ;
   RECT 0.0 112.86 272.84 114.57 ;
   RECT 0.0 114.57 272.84 116.28 ;
   RECT 0.0 116.28 272.84 117.99 ;
   RECT 0.0 117.99 272.84 119.7 ;
   RECT 0.0 119.7 272.84 121.41 ;
   RECT 0.0 121.41 272.84 123.12 ;
   RECT 0.0 123.12 272.84 124.83 ;
   RECT 0.0 124.83 296.02 126.54 ;
   RECT 0.0 126.54 296.02 128.25 ;
   RECT 0.0 128.25 296.02 129.96 ;
   RECT 0.0 129.96 296.02 131.67 ;
   RECT 0.0 131.67 296.02 133.38 ;
   RECT 0.0 133.38 296.02 135.09 ;
   RECT 0.0 135.09 296.02 136.8 ;
   RECT 0.0 136.8 296.02 138.51 ;
   RECT 0.0 138.51 296.02 140.22 ;
   RECT 0.0 140.22 296.02 141.93 ;
   RECT 0.0 141.93 296.02 143.64 ;
   RECT 0.0 143.64 296.02 145.35 ;
   RECT 0.0 145.35 296.02 147.06 ;
   RECT 0.0 147.06 296.02 148.77 ;
   RECT 0.0 148.77 296.02 150.48 ;
   RECT 0.0 150.48 296.02 152.19 ;
   RECT 0.0 152.19 296.02 153.9 ;
   RECT 0.0 153.9 272.84 155.61 ;
   RECT 0.0 155.61 272.84 157.32 ;
   RECT 0.0 157.32 272.84 159.03 ;
   RECT 0.0 159.03 272.84 160.74 ;
   RECT 0.0 160.74 272.84 162.45 ;
   RECT 0.0 162.45 272.84 164.16 ;
   RECT 0.0 164.16 272.84 165.87 ;
   RECT 0.0 165.87 272.84 167.58 ;
   RECT 0.0 167.58 272.84 169.29 ;
   RECT 0.0 169.29 272.84 171.0 ;
   RECT 0.0 171.0 272.84 172.71 ;
   RECT 0.0 172.71 272.84 174.42 ;
   RECT 0.0 174.42 272.84 176.13 ;
   RECT 0.0 176.13 272.84 177.84 ;
   RECT 0.0 177.84 272.84 179.55 ;
   RECT 0.0 179.55 272.84 181.26 ;
   RECT 0.0 181.26 272.84 182.97 ;
   RECT 0.0 182.97 272.84 184.68 ;
   RECT 0.0 184.68 272.84 186.39 ;
   RECT 0.0 186.39 272.84 188.1 ;
   RECT 0.0 188.1 272.84 189.81 ;
   RECT 0.0 189.81 272.84 191.52 ;
   RECT 0.0 191.52 272.84 193.23 ;
   RECT 0.0 193.23 272.84 194.94 ;
   RECT 0.0 194.94 272.84 196.65 ;
   RECT 0.0 196.65 272.84 198.36 ;
   RECT 0.0 198.36 272.84 200.07 ;
   RECT 0.0 200.07 272.84 201.78 ;
   RECT 0.0 201.78 272.84 203.49 ;
   RECT 0.0 203.49 272.84 205.2 ;
   RECT 0.0 205.2 272.84 206.91 ;
   RECT 0.0 206.91 272.84 208.62 ;
   RECT 0.0 208.62 272.84 210.33 ;
   RECT 0.0 210.33 272.84 212.04 ;
   RECT 0.0 212.04 272.84 213.75 ;
   RECT 0.0 213.75 272.84 215.46 ;
   RECT 0.0 215.46 272.84 217.17 ;
   RECT 0.0 217.17 272.84 218.88 ;
   RECT 0.0 218.88 272.84 220.59 ;
   RECT 0.0 220.59 272.84 222.3 ;
   RECT 0.0 222.3 272.84 224.01 ;
   RECT 0.0 224.01 272.84 225.72 ;
   RECT 0.0 225.72 272.84 227.43 ;
   RECT 0.0 227.43 272.84 229.14 ;
   RECT 0.0 229.14 272.84 230.85 ;
   RECT 0.0 230.85 272.84 232.56 ;
   RECT 0.0 232.56 272.84 234.27 ;
   RECT 0.0 234.27 272.84 235.98 ;
   RECT 0.0 235.98 272.84 237.69 ;
   RECT 0.0 237.69 272.84 239.4 ;
   RECT 0.0 239.4 272.84 241.11 ;
   RECT 0.0 241.11 272.84 242.82 ;
   RECT 0.0 242.82 272.84 244.53 ;
   RECT 0.0 244.53 272.84 246.24 ;
   RECT 0.0 246.24 272.84 247.95 ;
   RECT 0.0 247.95 272.84 249.66 ;
   RECT 0.0 249.66 272.84 251.37 ;
   RECT 0.0 251.37 272.84 253.08 ;
   RECT 0.0 253.08 272.84 254.79 ;
   RECT 0.0 254.79 272.84 256.5 ;
   RECT 0.0 256.5 272.84 258.21 ;
   RECT 0.0 258.21 272.84 259.92 ;
   RECT 0.0 259.92 272.84 261.63 ;
   RECT 0.0 261.63 272.84 263.34 ;
   RECT 0.0 263.34 272.84 265.05 ;
   RECT 0.0 265.05 272.84 266.76 ;
   RECT 0.0 266.76 272.84 268.47 ;
   RECT 0.0 268.47 272.84 270.18 ;
   RECT 0.0 270.18 272.84 271.89 ;
 END
END block_779x1431_153

MACRO block_546x675_104
 CLASS BLOCK ;
 FOREIGN block_546x675_104 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 207.48 BY 128.25 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 18.335 204.345 18.905 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 19.855 204.345 20.425 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 20.615 204.345 21.185 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 21.375 204.345 21.945 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 22.135 204.345 22.705 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 22.895 204.345 23.465 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 24.415 204.345 24.985 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 25.175 204.345 25.745 ;
  END
 END o7
 PIN o8
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 25.935 204.345 26.505 ;
  END
 END o8
 PIN o9
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 26.695 204.345 27.265 ;
  END
 END o9
 PIN o10
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 27.455 204.345 28.025 ;
  END
 END o10
 PIN o11
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 28.975 204.345 29.545 ;
  END
 END o11
 PIN o12
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 29.735 204.345 30.305 ;
  END
 END o12
 PIN o13
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 30.495 204.345 31.065 ;
  END
 END o13
 PIN o14
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 31.255 204.345 31.825 ;
  END
 END o14
 PIN o15
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 48.735 204.345 49.305 ;
  END
 END o15
 PIN o16
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 33.535 204.345 34.105 ;
  END
 END o16
 PIN o17
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 35.055 204.345 35.625 ;
  END
 END o17
 PIN o18
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 35.815 204.345 36.385 ;
  END
 END o18
 PIN o19
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 36.575 204.345 37.145 ;
  END
 END o19
 PIN o20
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 38.095 204.345 38.665 ;
  END
 END o20
 PIN o21
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 38.855 204.345 39.425 ;
  END
 END o21
 PIN o22
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 39.615 204.345 40.185 ;
  END
 END o22
 PIN o23
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 40.375 204.345 40.945 ;
  END
 END o23
 PIN o24
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 41.135 204.345 41.705 ;
  END
 END o24
 PIN o25
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 42.655 204.345 43.225 ;
  END
 END o25
 PIN o26
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 43.415 204.345 43.985 ;
  END
 END o26
 PIN o27
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 44.175 204.345 44.745 ;
  END
 END o27
 PIN o28
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 44.935 204.345 45.505 ;
  END
 END o28
 PIN o29
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 45.695 204.345 46.265 ;
  END
 END o29
 PIN o30
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 47.215 204.345 47.785 ;
  END
 END o30
 PIN o31
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 47.975 204.345 48.545 ;
  END
 END o31
 PIN o32
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 49.495 204.345 50.065 ;
  END
 END o32
 PIN o33
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 50.255 204.345 50.825 ;
  END
 END o33
 PIN o34
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 51.775 204.345 52.345 ;
  END
 END o34
 PIN o35
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 52.535 204.345 53.105 ;
  END
 END o35
 PIN o36
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 53.295 204.345 53.865 ;
  END
 END o36
 PIN o37
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 54.055 204.345 54.625 ;
  END
 END o37
 PIN o38
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 54.815 204.345 55.385 ;
  END
 END o38
 PIN o39
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 95.095 126.825 95.665 127.395 ;
  END
 END o39
 PIN o40
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 101.555 126.825 102.125 127.395 ;
  END
 END o40
 PIN o41
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 104.215 126.825 104.785 127.395 ;
  END
 END o41
 PIN o42
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 107.255 126.825 107.825 127.395 ;
  END
 END o42
 PIN o43
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 110.675 126.825 111.245 127.395 ;
  END
 END o43
 PIN o44
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 114.095 126.825 114.665 127.395 ;
  END
 END o44
 PIN o45
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.135 126.825 117.705 127.395 ;
  END
 END o45
 PIN o46
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 119.795 126.825 120.365 127.395 ;
  END
 END o46
 PIN o47
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 122.835 126.825 123.405 127.395 ;
  END
 END o47
 PIN o48
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 132.715 126.825 133.285 127.395 ;
  END
 END o48
 PIN o49
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 4.275 3.325 4.845 ;
  END
 END o49
 PIN o50
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 20.995 3.325 21.565 ;
  END
 END o50
 PIN o51
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 20.235 3.325 20.805 ;
  END
 END o51
 PIN o52
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 18.715 3.325 19.285 ;
  END
 END o52
 PIN o53
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 62.035 3.325 62.605 ;
  END
 END o53
 PIN o54
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 58.995 3.325 59.565 ;
  END
 END o54
 PIN o55
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 58.235 3.325 58.805 ;
  END
 END o55
 PIN o56
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 153.995 126.825 154.565 127.395 ;
  END
 END o56
 PIN o57
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 172.995 126.825 173.565 127.395 ;
  END
 END o57
 PIN o58
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 176.035 126.825 176.605 127.395 ;
  END
 END o58
 PIN o59
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 179.455 126.825 180.025 127.395 ;
  END
 END o59
 PIN o60
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 181.735 126.825 182.305 127.395 ;
  END
 END o60
 PIN o61
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 185.155 126.825 185.725 127.395 ;
  END
 END o61
 PIN o62
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 188.575 126.825 189.145 127.395 ;
  END
 END o62
 PIN o63
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 191.615 126.825 192.185 127.395 ;
  END
 END o63
 PIN o64
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 200.735 126.825 201.305 127.395 ;
  END
 END o64
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 82.935 126.825 83.505 127.395 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 70.395 126.825 70.965 127.395 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 85.975 126.825 86.545 127.395 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 41.895 126.825 42.465 127.395 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 44.935 126.825 45.505 127.395 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 48.355 126.825 48.925 127.395 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 51.775 126.825 52.345 127.395 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 54.815 126.825 55.385 127.395 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 57.475 126.825 58.045 127.395 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 60.515 126.825 61.085 127.395 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 63.935 126.825 64.505 127.395 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 88.635 126.825 89.205 127.395 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 73.055 126.825 73.625 127.395 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 91.675 126.825 92.245 127.395 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 98.515 126.825 99.085 127.395 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 126.825 130.245 127.395 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 150.955 126.825 151.525 127.395 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 197.315 126.825 197.885 127.395 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 56.335 204.345 56.905 ;
  END
 END i18
 PIN i19
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 57.095 204.345 57.665 ;
  END
 END i19
 PIN i20
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 57.855 204.345 58.425 ;
  END
 END i20
 PIN i21
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 58.615 204.345 59.185 ;
  END
 END i21
 PIN i22
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 59.375 204.345 59.945 ;
  END
 END i22
 PIN i23
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 60.895 204.345 61.465 ;
  END
 END i23
 PIN i24
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 61.655 204.345 62.225 ;
  END
 END i24
 PIN i25
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 63.175 204.345 63.745 ;
  END
 END i25
 PIN i26
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 63.935 204.345 64.505 ;
  END
 END i26
 PIN i27
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 65.455 204.345 66.025 ;
  END
 END i27
 PIN i28
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 66.215 204.345 66.785 ;
  END
 END i28
 PIN i29
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 66.975 204.345 67.545 ;
  END
 END i29
 PIN i30
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 67.735 204.345 68.305 ;
  END
 END i30
 PIN i31
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 68.495 204.345 69.065 ;
  END
 END i31
 PIN i32
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 74.955 3.325 75.525 ;
  END
 END i32
 PIN i33
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 75.715 3.325 76.285 ;
  END
 END i33
 PIN i34
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 76.475 3.325 77.045 ;
  END
 END i34
 PIN i35
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 77.235 3.325 77.805 ;
  END
 END i35
 PIN i36
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 77.995 3.325 78.565 ;
  END
 END i36
 PIN i37
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 79.515 3.325 80.085 ;
  END
 END i37
 PIN i38
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 80.275 3.325 80.845 ;
  END
 END i38
 OBS
  LAYER metal1 ;
   RECT 0 0 207.48 128.25 ;
  LAYER via1 ;
   RECT 0 0 207.48 128.25 ;
  LAYER metal2 ;
   RECT 0 0 207.48 128.25 ;
  LAYER via2 ;
   RECT 0 0 207.48 128.25 ;
  LAYER metal3 ;
   RECT 0 0 207.48 128.25 ;
  LAYER via3 ;
   RECT 0 0 207.48 128.25 ;
  LAYER metal4 ;
   RECT 0 0 207.48 128.25 ;
 END
END block_546x675_104

MACRO block_533x1044_173
 CLASS BLOCK ;
 FOREIGN block_533x1044_173 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 202.54 BY 198.36 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 4.275 176.225 4.845 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 8.455 176.225 9.025 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 63.365 176.225 63.935 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 67.545 176.225 68.115 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 71.535 176.225 72.105 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 75.715 176.225 76.285 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 79.705 176.225 80.275 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 83.885 176.225 84.455 ;
  END
 END o7
 PIN o8
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 112.005 176.225 112.575 ;
  END
 END o8
 PIN o9
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 116.185 176.225 116.755 ;
  END
 END o9
 PIN o10
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 120.175 176.225 120.745 ;
  END
 END o10
 PIN o11
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 124.355 176.225 124.925 ;
  END
 END o11
 PIN o12
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 12.445 176.225 13.015 ;
  END
 END o12
 PIN o13
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 128.345 176.225 128.915 ;
  END
 END o13
 PIN o14
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 132.525 176.225 133.095 ;
  END
 END o14
 PIN o15
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 136.515 176.225 137.085 ;
  END
 END o15
 PIN o16
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 140.695 176.225 141.265 ;
  END
 END o16
 PIN o17
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 162.925 176.225 163.495 ;
  END
 END o17
 PIN o18
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 167.105 176.225 167.675 ;
  END
 END o18
 PIN o19
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 171.095 176.225 171.665 ;
  END
 END o19
 PIN o20
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 175.275 176.225 175.845 ;
  END
 END o20
 PIN o21
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 179.265 176.225 179.835 ;
  END
 END o21
 PIN o22
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 183.445 176.225 184.015 ;
  END
 END o22
 PIN o23
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 16.625 176.225 17.195 ;
  END
 END o23
 PIN o24
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 187.435 176.225 188.005 ;
  END
 END o24
 PIN o25
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 191.615 176.225 192.185 ;
  END
 END o25
 PIN o26
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 20.615 176.225 21.185 ;
  END
 END o26
 PIN o27
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 24.795 176.225 25.365 ;
  END
 END o27
 PIN o28
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 28.785 176.225 29.355 ;
  END
 END o28
 PIN o29
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 32.965 176.225 33.535 ;
  END
 END o29
 PIN o30
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 55.195 176.225 55.765 ;
  END
 END o30
 PIN o31
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 59.375 176.225 59.945 ;
  END
 END o31
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.835 86.735 199.405 87.305 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.835 103.835 199.405 104.405 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.835 92.055 199.405 92.625 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.075 87.115 198.645 87.685 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.075 86.355 198.645 86.925 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.835 85.975 199.405 86.545 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.835 95.665 199.405 96.235 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.835 108.775 199.405 109.345 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.075 103.455 198.645 104.025 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.835 103.075 199.405 103.645 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.835 105.165 199.405 105.735 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.835 107.635 199.405 108.205 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.075 109.155 198.645 109.725 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 188.955 85.595 189.525 86.165 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 188.955 98.895 189.525 99.465 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 2.565 176.225 3.135 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 6.745 176.225 7.315 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 61.655 176.225 62.225 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 65.835 176.225 66.405 ;
  END
 END i18
 PIN i19
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 69.825 176.225 70.395 ;
  END
 END i19
 PIN i20
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 74.005 176.225 74.575 ;
  END
 END i20
 PIN i21
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 77.995 176.225 78.565 ;
  END
 END i21
 PIN i22
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 82.175 176.225 82.745 ;
  END
 END i22
 PIN i23
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 113.715 176.225 114.285 ;
  END
 END i23
 PIN i24
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 117.895 176.225 118.465 ;
  END
 END i24
 PIN i25
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 121.885 176.225 122.455 ;
  END
 END i25
 PIN i26
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 126.065 176.225 126.635 ;
  END
 END i26
 PIN i27
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 10.735 176.225 11.305 ;
  END
 END i27
 PIN i28
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 130.055 176.225 130.625 ;
  END
 END i28
 PIN i29
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 134.235 176.225 134.805 ;
  END
 END i29
 PIN i30
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 138.225 176.225 138.795 ;
  END
 END i30
 PIN i31
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 142.405 176.225 142.975 ;
  END
 END i31
 PIN i32
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 164.635 176.225 165.205 ;
  END
 END i32
 PIN i33
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 168.815 176.225 169.385 ;
  END
 END i33
 PIN i34
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 172.805 176.225 173.375 ;
  END
 END i34
 PIN i35
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 176.985 176.225 177.555 ;
  END
 END i35
 PIN i36
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 180.975 176.225 181.545 ;
  END
 END i36
 PIN i37
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 185.155 176.225 185.725 ;
  END
 END i37
 PIN i38
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 14.915 176.225 15.485 ;
  END
 END i38
 PIN i39
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 189.145 176.225 189.715 ;
  END
 END i39
 PIN i40
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 193.325 176.225 193.895 ;
  END
 END i40
 PIN i41
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 18.905 176.225 19.475 ;
  END
 END i41
 PIN i42
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 23.085 176.225 23.655 ;
  END
 END i42
 PIN i43
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 27.075 176.225 27.645 ;
  END
 END i43
 PIN i44
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 31.255 176.225 31.825 ;
  END
 END i44
 PIN i45
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 53.485 176.225 54.055 ;
  END
 END i45
 PIN i46
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 57.665 176.225 58.235 ;
  END
 END i46
 PIN i47
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 9.025 175.465 9.595 ;
  END
 END i47
 PIN i48
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 13.015 175.465 13.585 ;
  END
 END i48
 PIN i49
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 17.195 175.465 17.765 ;
  END
 END i49
 PIN i50
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 76.285 175.465 76.855 ;
  END
 END i50
 PIN i51
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 80.275 175.465 80.845 ;
  END
 END i51
 PIN i52
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 84.455 175.465 85.025 ;
  END
 END i52
 PIN i53
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 119.605 175.465 120.175 ;
  END
 END i53
 PIN i54
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 115.615 175.465 116.185 ;
  END
 END i54
 PIN i55
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 111.435 175.465 112.005 ;
  END
 END i55
 PIN i56
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 186.865 175.465 187.435 ;
  END
 END i56
 PIN i57
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 182.875 175.465 183.445 ;
  END
 END i57
 PIN i58
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 178.695 175.465 179.265 ;
  END
 END i58
 PIN i59
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 4.845 175.465 5.415 ;
  END
 END i59
 PIN i60
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 72.105 175.465 72.675 ;
  END
 END i60
 PIN i61
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 123.785 175.465 124.355 ;
  END
 END i61
 PIN i62
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 191.045 175.465 191.615 ;
  END
 END i62
 PIN i63
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 184.015 85.595 184.585 86.165 ;
  END
 END i63
 PIN i64
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 184.015 98.895 184.585 99.465 ;
  END
 END i64
 PIN i65
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 3.135 175.465 3.705 ;
  END
 END i65
 PIN i66
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 7.315 175.465 7.885 ;
  END
 END i66
 PIN i67
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 62.225 175.465 62.795 ;
  END
 END i67
 PIN i68
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 66.405 175.465 66.975 ;
  END
 END i68
 PIN i69
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 70.395 175.465 70.965 ;
  END
 END i69
 PIN i70
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 74.575 175.465 75.145 ;
  END
 END i70
 PIN i71
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 78.565 175.465 79.135 ;
  END
 END i71
 PIN i72
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 82.745 175.465 83.315 ;
  END
 END i72
 PIN i73
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 113.145 175.465 113.715 ;
  END
 END i73
 PIN i74
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 117.325 175.465 117.895 ;
  END
 END i74
 PIN i75
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 121.315 175.465 121.885 ;
  END
 END i75
 PIN i76
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 125.495 175.465 126.065 ;
  END
 END i76
 PIN i77
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 11.305 175.465 11.875 ;
  END
 END i77
 PIN i78
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 129.485 175.465 130.055 ;
  END
 END i78
 PIN i79
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 133.665 175.465 134.235 ;
  END
 END i79
 PIN i80
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 137.655 175.465 138.225 ;
  END
 END i80
 PIN i81
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 141.835 175.465 142.405 ;
  END
 END i81
 PIN i82
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 164.065 175.465 164.635 ;
  END
 END i82
 PIN i83
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 168.245 175.465 168.815 ;
  END
 END i83
 PIN i84
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 172.235 175.465 172.805 ;
  END
 END i84
 PIN i85
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 176.415 175.465 176.985 ;
  END
 END i85
 PIN i86
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 180.405 175.465 180.975 ;
  END
 END i86
 PIN i87
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 184.585 175.465 185.155 ;
  END
 END i87
 PIN i88
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 15.485 175.465 16.055 ;
  END
 END i88
 PIN i89
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 188.575 175.465 189.145 ;
  END
 END i89
 PIN i90
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 192.755 175.465 193.325 ;
  END
 END i90
 PIN i91
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 19.475 175.465 20.045 ;
  END
 END i91
 PIN i92
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 23.655 175.465 24.225 ;
  END
 END i92
 PIN i93
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 27.645 175.465 28.215 ;
  END
 END i93
 PIN i94
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 31.825 175.465 32.395 ;
  END
 END i94
 PIN i95
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 54.055 175.465 54.625 ;
  END
 END i95
 PIN i96
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 58.235 175.465 58.805 ;
  END
 END i96
 PIN i97
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.835 93.195 199.405 93.765 ;
  END
 END i97
 PIN i98
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.075 93.575 198.645 94.145 ;
  END
 END i98
 PIN i99
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 3.705 174.705 4.275 ;
  END
 END i99
 PIN i100
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 7.885 174.705 8.455 ;
  END
 END i100
 PIN i101
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 62.795 174.705 63.365 ;
  END
 END i101
 PIN i102
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 66.975 174.705 67.545 ;
  END
 END i102
 PIN i103
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 70.965 174.705 71.535 ;
  END
 END i103
 PIN i104
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 75.145 174.705 75.715 ;
  END
 END i104
 PIN i105
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 79.135 174.705 79.705 ;
  END
 END i105
 PIN i106
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 83.315 174.705 83.885 ;
  END
 END i106
 PIN i107
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 112.575 174.705 113.145 ;
  END
 END i107
 PIN i108
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 116.755 174.705 117.325 ;
  END
 END i108
 PIN i109
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 120.745 174.705 121.315 ;
  END
 END i109
 PIN i110
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 124.925 174.705 125.495 ;
  END
 END i110
 PIN i111
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 11.875 174.705 12.445 ;
  END
 END i111
 PIN i112
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 128.915 174.705 129.485 ;
  END
 END i112
 PIN i113
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 133.095 174.705 133.665 ;
  END
 END i113
 PIN i114
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 137.085 174.705 137.655 ;
  END
 END i114
 PIN i115
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 141.265 174.705 141.835 ;
  END
 END i115
 PIN i116
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 163.495 174.705 164.065 ;
  END
 END i116
 PIN i117
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 167.675 174.705 168.245 ;
  END
 END i117
 PIN i118
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 171.665 174.705 172.235 ;
  END
 END i118
 PIN i119
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 175.845 174.705 176.415 ;
  END
 END i119
 PIN i120
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 179.835 174.705 180.405 ;
  END
 END i120
 PIN i121
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 184.015 174.705 184.585 ;
  END
 END i121
 PIN i122
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 16.055 174.705 16.625 ;
  END
 END i122
 PIN i123
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 188.005 174.705 188.575 ;
  END
 END i123
 PIN i124
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 192.185 174.705 192.755 ;
  END
 END i124
 PIN i125
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 20.045 174.705 20.615 ;
  END
 END i125
 PIN i126
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 24.225 174.705 24.795 ;
  END
 END i126
 PIN i127
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 28.215 174.705 28.785 ;
  END
 END i127
 PIN i128
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 32.395 174.705 32.965 ;
  END
 END i128
 PIN i129
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 54.625 174.705 55.195 ;
  END
 END i129
 PIN i130
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 58.805 174.705 59.375 ;
  END
 END i130
 PIN i131
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 197.695 85.595 198.265 86.165 ;
  END
 END i131
 PIN i132
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 196.555 85.595 197.125 86.165 ;
  END
 END i132
 PIN i133
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 195.035 85.595 195.605 86.165 ;
  END
 END i133
 PIN i134
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 193.135 85.595 193.705 86.165 ;
  END
 END i134
 PIN i135
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 191.995 85.595 192.565 86.165 ;
  END
 END i135
 PIN i136
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 197.695 98.895 198.265 99.465 ;
  END
 END i136
 PIN i137
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 196.555 98.895 197.125 99.465 ;
  END
 END i137
 PIN i138
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 195.035 98.895 195.605 99.465 ;
  END
 END i138
 PIN i139
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 193.135 98.895 193.705 99.465 ;
  END
 END i139
 PIN i140
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 191.995 98.895 192.565 99.465 ;
  END
 END i140
 OBS
  LAYER metal1 ;
   RECT 0.0 0.0 179.36 1.71 ;
   RECT 0.0 1.71 179.36 3.42 ;
   RECT 0.0 3.42 179.36 5.13 ;
   RECT 0.0 5.13 179.36 6.84 ;
   RECT 0.0 6.84 179.36 8.55 ;
   RECT 0.0 8.55 179.36 10.26 ;
   RECT 0.0 10.26 179.36 11.97 ;
   RECT 0.0 11.97 179.36 13.68 ;
   RECT 0.0 13.68 179.36 15.39 ;
   RECT 0.0 15.39 179.36 17.1 ;
   RECT 0.0 17.1 179.36 18.81 ;
   RECT 0.0 18.81 179.36 20.52 ;
   RECT 0.0 20.52 179.36 22.23 ;
   RECT 0.0 22.23 179.36 23.94 ;
   RECT 0.0 23.94 179.36 25.65 ;
   RECT 0.0 25.65 179.36 27.36 ;
   RECT 0.0 27.36 179.36 29.07 ;
   RECT 0.0 29.07 179.36 30.78 ;
   RECT 0.0 30.78 179.36 32.49 ;
   RECT 0.0 32.49 179.36 34.2 ;
   RECT 0.0 34.2 179.36 35.91 ;
   RECT 0.0 35.91 179.36 37.62 ;
   RECT 0.0 37.62 179.36 39.33 ;
   RECT 0.0 39.33 179.36 41.04 ;
   RECT 0.0 41.04 179.36 42.75 ;
   RECT 0.0 42.75 179.36 44.46 ;
   RECT 0.0 44.46 179.36 46.17 ;
   RECT 0.0 46.17 179.36 47.88 ;
   RECT 0.0 47.88 179.36 49.59 ;
   RECT 0.0 49.59 179.36 51.3 ;
   RECT 0.0 51.3 179.36 53.01 ;
   RECT 0.0 53.01 179.36 54.72 ;
   RECT 0.0 54.72 179.36 56.43 ;
   RECT 0.0 56.43 179.36 58.14 ;
   RECT 0.0 58.14 179.36 59.85 ;
   RECT 0.0 59.85 179.36 61.56 ;
   RECT 0.0 61.56 179.36 63.27 ;
   RECT 0.0 63.27 179.36 64.98 ;
   RECT 0.0 64.98 179.36 66.69 ;
   RECT 0.0 66.69 179.36 68.4 ;
   RECT 0.0 68.4 179.36 70.11 ;
   RECT 0.0 70.11 179.36 71.82 ;
   RECT 0.0 71.82 179.36 73.53 ;
   RECT 0.0 73.53 179.36 75.24 ;
   RECT 0.0 75.24 179.36 76.95 ;
   RECT 0.0 76.95 179.36 78.66 ;
   RECT 0.0 78.66 179.36 80.37 ;
   RECT 0.0 80.37 179.36 82.08 ;
   RECT 0.0 82.08 179.36 83.79 ;
   RECT 0.0 83.79 202.54 85.5 ;
   RECT 0.0 85.5 202.54 87.21 ;
   RECT 0.0 87.21 202.54 88.92 ;
   RECT 0.0 88.92 202.54 90.63 ;
   RECT 0.0 90.63 202.54 92.34 ;
   RECT 0.0 92.34 202.54 94.05 ;
   RECT 0.0 94.05 202.54 95.76 ;
   RECT 0.0 95.76 202.54 97.47 ;
   RECT 0.0 97.47 202.54 99.18 ;
   RECT 0.0 99.18 202.54 100.89 ;
   RECT 0.0 100.89 202.54 102.6 ;
   RECT 0.0 102.6 202.54 104.31 ;
   RECT 0.0 104.31 202.54 106.02 ;
   RECT 0.0 106.02 202.54 107.73 ;
   RECT 0.0 107.73 202.54 109.44 ;
   RECT 0.0 109.44 202.54 111.15 ;
   RECT 0.0 111.15 202.54 112.86 ;
   RECT 0.0 112.86 179.36 114.57 ;
   RECT 0.0 114.57 179.36 116.28 ;
   RECT 0.0 116.28 179.36 117.99 ;
   RECT 0.0 117.99 179.36 119.7 ;
   RECT 0.0 119.7 179.36 121.41 ;
   RECT 0.0 121.41 179.36 123.12 ;
   RECT 0.0 123.12 179.36 124.83 ;
   RECT 0.0 124.83 179.36 126.54 ;
   RECT 0.0 126.54 179.36 128.25 ;
   RECT 0.0 128.25 179.36 129.96 ;
   RECT 0.0 129.96 179.36 131.67 ;
   RECT 0.0 131.67 179.36 133.38 ;
   RECT 0.0 133.38 179.36 135.09 ;
   RECT 0.0 135.09 179.36 136.8 ;
   RECT 0.0 136.8 179.36 138.51 ;
   RECT 0.0 138.51 179.36 140.22 ;
   RECT 0.0 140.22 179.36 141.93 ;
   RECT 0.0 141.93 179.36 143.64 ;
   RECT 0.0 143.64 179.36 145.35 ;
   RECT 0.0 145.35 179.36 147.06 ;
   RECT 0.0 147.06 179.36 148.77 ;
   RECT 0.0 148.77 179.36 150.48 ;
   RECT 0.0 150.48 179.36 152.19 ;
   RECT 0.0 152.19 179.36 153.9 ;
   RECT 0.0 153.9 179.36 155.61 ;
   RECT 0.0 155.61 179.36 157.32 ;
   RECT 0.0 157.32 179.36 159.03 ;
   RECT 0.0 159.03 179.36 160.74 ;
   RECT 0.0 160.74 179.36 162.45 ;
   RECT 0.0 162.45 179.36 164.16 ;
   RECT 0.0 164.16 179.36 165.87 ;
   RECT 0.0 165.87 179.36 167.58 ;
   RECT 0.0 167.58 179.36 169.29 ;
   RECT 0.0 169.29 179.36 171.0 ;
   RECT 0.0 171.0 179.36 172.71 ;
   RECT 0.0 172.71 179.36 174.42 ;
   RECT 0.0 174.42 179.36 176.13 ;
   RECT 0.0 176.13 179.36 177.84 ;
   RECT 0.0 177.84 179.36 179.55 ;
   RECT 0.0 179.55 179.36 181.26 ;
   RECT 0.0 181.26 179.36 182.97 ;
   RECT 0.0 182.97 179.36 184.68 ;
   RECT 0.0 184.68 179.36 186.39 ;
   RECT 0.0 186.39 179.36 188.1 ;
   RECT 0.0 188.1 179.36 189.81 ;
   RECT 0.0 189.81 179.36 191.52 ;
   RECT 0.0 191.52 179.36 193.23 ;
   RECT 0.0 193.23 179.36 194.94 ;
   RECT 0.0 194.94 179.36 196.65 ;
   RECT 0.0 196.65 179.36 198.36 ;
  LAYER via1 ;
   RECT 0.0 0.0 179.36 1.71 ;
   RECT 0.0 1.71 179.36 3.42 ;
   RECT 0.0 3.42 179.36 5.13 ;
   RECT 0.0 5.13 179.36 6.84 ;
   RECT 0.0 6.84 179.36 8.55 ;
   RECT 0.0 8.55 179.36 10.26 ;
   RECT 0.0 10.26 179.36 11.97 ;
   RECT 0.0 11.97 179.36 13.68 ;
   RECT 0.0 13.68 179.36 15.39 ;
   RECT 0.0 15.39 179.36 17.1 ;
   RECT 0.0 17.1 179.36 18.81 ;
   RECT 0.0 18.81 179.36 20.52 ;
   RECT 0.0 20.52 179.36 22.23 ;
   RECT 0.0 22.23 179.36 23.94 ;
   RECT 0.0 23.94 179.36 25.65 ;
   RECT 0.0 25.65 179.36 27.36 ;
   RECT 0.0 27.36 179.36 29.07 ;
   RECT 0.0 29.07 179.36 30.78 ;
   RECT 0.0 30.78 179.36 32.49 ;
   RECT 0.0 32.49 179.36 34.2 ;
   RECT 0.0 34.2 179.36 35.91 ;
   RECT 0.0 35.91 179.36 37.62 ;
   RECT 0.0 37.62 179.36 39.33 ;
   RECT 0.0 39.33 179.36 41.04 ;
   RECT 0.0 41.04 179.36 42.75 ;
   RECT 0.0 42.75 179.36 44.46 ;
   RECT 0.0 44.46 179.36 46.17 ;
   RECT 0.0 46.17 179.36 47.88 ;
   RECT 0.0 47.88 179.36 49.59 ;
   RECT 0.0 49.59 179.36 51.3 ;
   RECT 0.0 51.3 179.36 53.01 ;
   RECT 0.0 53.01 179.36 54.72 ;
   RECT 0.0 54.72 179.36 56.43 ;
   RECT 0.0 56.43 179.36 58.14 ;
   RECT 0.0 58.14 179.36 59.85 ;
   RECT 0.0 59.85 179.36 61.56 ;
   RECT 0.0 61.56 179.36 63.27 ;
   RECT 0.0 63.27 179.36 64.98 ;
   RECT 0.0 64.98 179.36 66.69 ;
   RECT 0.0 66.69 179.36 68.4 ;
   RECT 0.0 68.4 179.36 70.11 ;
   RECT 0.0 70.11 179.36 71.82 ;
   RECT 0.0 71.82 179.36 73.53 ;
   RECT 0.0 73.53 179.36 75.24 ;
   RECT 0.0 75.24 179.36 76.95 ;
   RECT 0.0 76.95 179.36 78.66 ;
   RECT 0.0 78.66 179.36 80.37 ;
   RECT 0.0 80.37 179.36 82.08 ;
   RECT 0.0 82.08 179.36 83.79 ;
   RECT 0.0 83.79 202.54 85.5 ;
   RECT 0.0 85.5 202.54 87.21 ;
   RECT 0.0 87.21 202.54 88.92 ;
   RECT 0.0 88.92 202.54 90.63 ;
   RECT 0.0 90.63 202.54 92.34 ;
   RECT 0.0 92.34 202.54 94.05 ;
   RECT 0.0 94.05 202.54 95.76 ;
   RECT 0.0 95.76 202.54 97.47 ;
   RECT 0.0 97.47 202.54 99.18 ;
   RECT 0.0 99.18 202.54 100.89 ;
   RECT 0.0 100.89 202.54 102.6 ;
   RECT 0.0 102.6 202.54 104.31 ;
   RECT 0.0 104.31 202.54 106.02 ;
   RECT 0.0 106.02 202.54 107.73 ;
   RECT 0.0 107.73 202.54 109.44 ;
   RECT 0.0 109.44 202.54 111.15 ;
   RECT 0.0 111.15 202.54 112.86 ;
   RECT 0.0 112.86 179.36 114.57 ;
   RECT 0.0 114.57 179.36 116.28 ;
   RECT 0.0 116.28 179.36 117.99 ;
   RECT 0.0 117.99 179.36 119.7 ;
   RECT 0.0 119.7 179.36 121.41 ;
   RECT 0.0 121.41 179.36 123.12 ;
   RECT 0.0 123.12 179.36 124.83 ;
   RECT 0.0 124.83 179.36 126.54 ;
   RECT 0.0 126.54 179.36 128.25 ;
   RECT 0.0 128.25 179.36 129.96 ;
   RECT 0.0 129.96 179.36 131.67 ;
   RECT 0.0 131.67 179.36 133.38 ;
   RECT 0.0 133.38 179.36 135.09 ;
   RECT 0.0 135.09 179.36 136.8 ;
   RECT 0.0 136.8 179.36 138.51 ;
   RECT 0.0 138.51 179.36 140.22 ;
   RECT 0.0 140.22 179.36 141.93 ;
   RECT 0.0 141.93 179.36 143.64 ;
   RECT 0.0 143.64 179.36 145.35 ;
   RECT 0.0 145.35 179.36 147.06 ;
   RECT 0.0 147.06 179.36 148.77 ;
   RECT 0.0 148.77 179.36 150.48 ;
   RECT 0.0 150.48 179.36 152.19 ;
   RECT 0.0 152.19 179.36 153.9 ;
   RECT 0.0 153.9 179.36 155.61 ;
   RECT 0.0 155.61 179.36 157.32 ;
   RECT 0.0 157.32 179.36 159.03 ;
   RECT 0.0 159.03 179.36 160.74 ;
   RECT 0.0 160.74 179.36 162.45 ;
   RECT 0.0 162.45 179.36 164.16 ;
   RECT 0.0 164.16 179.36 165.87 ;
   RECT 0.0 165.87 179.36 167.58 ;
   RECT 0.0 167.58 179.36 169.29 ;
   RECT 0.0 169.29 179.36 171.0 ;
   RECT 0.0 171.0 179.36 172.71 ;
   RECT 0.0 172.71 179.36 174.42 ;
   RECT 0.0 174.42 179.36 176.13 ;
   RECT 0.0 176.13 179.36 177.84 ;
   RECT 0.0 177.84 179.36 179.55 ;
   RECT 0.0 179.55 179.36 181.26 ;
   RECT 0.0 181.26 179.36 182.97 ;
   RECT 0.0 182.97 179.36 184.68 ;
   RECT 0.0 184.68 179.36 186.39 ;
   RECT 0.0 186.39 179.36 188.1 ;
   RECT 0.0 188.1 179.36 189.81 ;
   RECT 0.0 189.81 179.36 191.52 ;
   RECT 0.0 191.52 179.36 193.23 ;
   RECT 0.0 193.23 179.36 194.94 ;
   RECT 0.0 194.94 179.36 196.65 ;
   RECT 0.0 196.65 179.36 198.36 ;
  LAYER metal2 ;
   RECT 0.0 0.0 179.36 1.71 ;
   RECT 0.0 1.71 179.36 3.42 ;
   RECT 0.0 3.42 179.36 5.13 ;
   RECT 0.0 5.13 179.36 6.84 ;
   RECT 0.0 6.84 179.36 8.55 ;
   RECT 0.0 8.55 179.36 10.26 ;
   RECT 0.0 10.26 179.36 11.97 ;
   RECT 0.0 11.97 179.36 13.68 ;
   RECT 0.0 13.68 179.36 15.39 ;
   RECT 0.0 15.39 179.36 17.1 ;
   RECT 0.0 17.1 179.36 18.81 ;
   RECT 0.0 18.81 179.36 20.52 ;
   RECT 0.0 20.52 179.36 22.23 ;
   RECT 0.0 22.23 179.36 23.94 ;
   RECT 0.0 23.94 179.36 25.65 ;
   RECT 0.0 25.65 179.36 27.36 ;
   RECT 0.0 27.36 179.36 29.07 ;
   RECT 0.0 29.07 179.36 30.78 ;
   RECT 0.0 30.78 179.36 32.49 ;
   RECT 0.0 32.49 179.36 34.2 ;
   RECT 0.0 34.2 179.36 35.91 ;
   RECT 0.0 35.91 179.36 37.62 ;
   RECT 0.0 37.62 179.36 39.33 ;
   RECT 0.0 39.33 179.36 41.04 ;
   RECT 0.0 41.04 179.36 42.75 ;
   RECT 0.0 42.75 179.36 44.46 ;
   RECT 0.0 44.46 179.36 46.17 ;
   RECT 0.0 46.17 179.36 47.88 ;
   RECT 0.0 47.88 179.36 49.59 ;
   RECT 0.0 49.59 179.36 51.3 ;
   RECT 0.0 51.3 179.36 53.01 ;
   RECT 0.0 53.01 179.36 54.72 ;
   RECT 0.0 54.72 179.36 56.43 ;
   RECT 0.0 56.43 179.36 58.14 ;
   RECT 0.0 58.14 179.36 59.85 ;
   RECT 0.0 59.85 179.36 61.56 ;
   RECT 0.0 61.56 179.36 63.27 ;
   RECT 0.0 63.27 179.36 64.98 ;
   RECT 0.0 64.98 179.36 66.69 ;
   RECT 0.0 66.69 179.36 68.4 ;
   RECT 0.0 68.4 179.36 70.11 ;
   RECT 0.0 70.11 179.36 71.82 ;
   RECT 0.0 71.82 179.36 73.53 ;
   RECT 0.0 73.53 179.36 75.24 ;
   RECT 0.0 75.24 179.36 76.95 ;
   RECT 0.0 76.95 179.36 78.66 ;
   RECT 0.0 78.66 179.36 80.37 ;
   RECT 0.0 80.37 179.36 82.08 ;
   RECT 0.0 82.08 179.36 83.79 ;
   RECT 0.0 83.79 202.54 85.5 ;
   RECT 0.0 85.5 202.54 87.21 ;
   RECT 0.0 87.21 202.54 88.92 ;
   RECT 0.0 88.92 202.54 90.63 ;
   RECT 0.0 90.63 202.54 92.34 ;
   RECT 0.0 92.34 202.54 94.05 ;
   RECT 0.0 94.05 202.54 95.76 ;
   RECT 0.0 95.76 202.54 97.47 ;
   RECT 0.0 97.47 202.54 99.18 ;
   RECT 0.0 99.18 202.54 100.89 ;
   RECT 0.0 100.89 202.54 102.6 ;
   RECT 0.0 102.6 202.54 104.31 ;
   RECT 0.0 104.31 202.54 106.02 ;
   RECT 0.0 106.02 202.54 107.73 ;
   RECT 0.0 107.73 202.54 109.44 ;
   RECT 0.0 109.44 202.54 111.15 ;
   RECT 0.0 111.15 202.54 112.86 ;
   RECT 0.0 112.86 179.36 114.57 ;
   RECT 0.0 114.57 179.36 116.28 ;
   RECT 0.0 116.28 179.36 117.99 ;
   RECT 0.0 117.99 179.36 119.7 ;
   RECT 0.0 119.7 179.36 121.41 ;
   RECT 0.0 121.41 179.36 123.12 ;
   RECT 0.0 123.12 179.36 124.83 ;
   RECT 0.0 124.83 179.36 126.54 ;
   RECT 0.0 126.54 179.36 128.25 ;
   RECT 0.0 128.25 179.36 129.96 ;
   RECT 0.0 129.96 179.36 131.67 ;
   RECT 0.0 131.67 179.36 133.38 ;
   RECT 0.0 133.38 179.36 135.09 ;
   RECT 0.0 135.09 179.36 136.8 ;
   RECT 0.0 136.8 179.36 138.51 ;
   RECT 0.0 138.51 179.36 140.22 ;
   RECT 0.0 140.22 179.36 141.93 ;
   RECT 0.0 141.93 179.36 143.64 ;
   RECT 0.0 143.64 179.36 145.35 ;
   RECT 0.0 145.35 179.36 147.06 ;
   RECT 0.0 147.06 179.36 148.77 ;
   RECT 0.0 148.77 179.36 150.48 ;
   RECT 0.0 150.48 179.36 152.19 ;
   RECT 0.0 152.19 179.36 153.9 ;
   RECT 0.0 153.9 179.36 155.61 ;
   RECT 0.0 155.61 179.36 157.32 ;
   RECT 0.0 157.32 179.36 159.03 ;
   RECT 0.0 159.03 179.36 160.74 ;
   RECT 0.0 160.74 179.36 162.45 ;
   RECT 0.0 162.45 179.36 164.16 ;
   RECT 0.0 164.16 179.36 165.87 ;
   RECT 0.0 165.87 179.36 167.58 ;
   RECT 0.0 167.58 179.36 169.29 ;
   RECT 0.0 169.29 179.36 171.0 ;
   RECT 0.0 171.0 179.36 172.71 ;
   RECT 0.0 172.71 179.36 174.42 ;
   RECT 0.0 174.42 179.36 176.13 ;
   RECT 0.0 176.13 179.36 177.84 ;
   RECT 0.0 177.84 179.36 179.55 ;
   RECT 0.0 179.55 179.36 181.26 ;
   RECT 0.0 181.26 179.36 182.97 ;
   RECT 0.0 182.97 179.36 184.68 ;
   RECT 0.0 184.68 179.36 186.39 ;
   RECT 0.0 186.39 179.36 188.1 ;
   RECT 0.0 188.1 179.36 189.81 ;
   RECT 0.0 189.81 179.36 191.52 ;
   RECT 0.0 191.52 179.36 193.23 ;
   RECT 0.0 193.23 179.36 194.94 ;
   RECT 0.0 194.94 179.36 196.65 ;
   RECT 0.0 196.65 179.36 198.36 ;
  LAYER via2 ;
   RECT 0.0 0.0 179.36 1.71 ;
   RECT 0.0 1.71 179.36 3.42 ;
   RECT 0.0 3.42 179.36 5.13 ;
   RECT 0.0 5.13 179.36 6.84 ;
   RECT 0.0 6.84 179.36 8.55 ;
   RECT 0.0 8.55 179.36 10.26 ;
   RECT 0.0 10.26 179.36 11.97 ;
   RECT 0.0 11.97 179.36 13.68 ;
   RECT 0.0 13.68 179.36 15.39 ;
   RECT 0.0 15.39 179.36 17.1 ;
   RECT 0.0 17.1 179.36 18.81 ;
   RECT 0.0 18.81 179.36 20.52 ;
   RECT 0.0 20.52 179.36 22.23 ;
   RECT 0.0 22.23 179.36 23.94 ;
   RECT 0.0 23.94 179.36 25.65 ;
   RECT 0.0 25.65 179.36 27.36 ;
   RECT 0.0 27.36 179.36 29.07 ;
   RECT 0.0 29.07 179.36 30.78 ;
   RECT 0.0 30.78 179.36 32.49 ;
   RECT 0.0 32.49 179.36 34.2 ;
   RECT 0.0 34.2 179.36 35.91 ;
   RECT 0.0 35.91 179.36 37.62 ;
   RECT 0.0 37.62 179.36 39.33 ;
   RECT 0.0 39.33 179.36 41.04 ;
   RECT 0.0 41.04 179.36 42.75 ;
   RECT 0.0 42.75 179.36 44.46 ;
   RECT 0.0 44.46 179.36 46.17 ;
   RECT 0.0 46.17 179.36 47.88 ;
   RECT 0.0 47.88 179.36 49.59 ;
   RECT 0.0 49.59 179.36 51.3 ;
   RECT 0.0 51.3 179.36 53.01 ;
   RECT 0.0 53.01 179.36 54.72 ;
   RECT 0.0 54.72 179.36 56.43 ;
   RECT 0.0 56.43 179.36 58.14 ;
   RECT 0.0 58.14 179.36 59.85 ;
   RECT 0.0 59.85 179.36 61.56 ;
   RECT 0.0 61.56 179.36 63.27 ;
   RECT 0.0 63.27 179.36 64.98 ;
   RECT 0.0 64.98 179.36 66.69 ;
   RECT 0.0 66.69 179.36 68.4 ;
   RECT 0.0 68.4 179.36 70.11 ;
   RECT 0.0 70.11 179.36 71.82 ;
   RECT 0.0 71.82 179.36 73.53 ;
   RECT 0.0 73.53 179.36 75.24 ;
   RECT 0.0 75.24 179.36 76.95 ;
   RECT 0.0 76.95 179.36 78.66 ;
   RECT 0.0 78.66 179.36 80.37 ;
   RECT 0.0 80.37 179.36 82.08 ;
   RECT 0.0 82.08 179.36 83.79 ;
   RECT 0.0 83.79 202.54 85.5 ;
   RECT 0.0 85.5 202.54 87.21 ;
   RECT 0.0 87.21 202.54 88.92 ;
   RECT 0.0 88.92 202.54 90.63 ;
   RECT 0.0 90.63 202.54 92.34 ;
   RECT 0.0 92.34 202.54 94.05 ;
   RECT 0.0 94.05 202.54 95.76 ;
   RECT 0.0 95.76 202.54 97.47 ;
   RECT 0.0 97.47 202.54 99.18 ;
   RECT 0.0 99.18 202.54 100.89 ;
   RECT 0.0 100.89 202.54 102.6 ;
   RECT 0.0 102.6 202.54 104.31 ;
   RECT 0.0 104.31 202.54 106.02 ;
   RECT 0.0 106.02 202.54 107.73 ;
   RECT 0.0 107.73 202.54 109.44 ;
   RECT 0.0 109.44 202.54 111.15 ;
   RECT 0.0 111.15 202.54 112.86 ;
   RECT 0.0 112.86 179.36 114.57 ;
   RECT 0.0 114.57 179.36 116.28 ;
   RECT 0.0 116.28 179.36 117.99 ;
   RECT 0.0 117.99 179.36 119.7 ;
   RECT 0.0 119.7 179.36 121.41 ;
   RECT 0.0 121.41 179.36 123.12 ;
   RECT 0.0 123.12 179.36 124.83 ;
   RECT 0.0 124.83 179.36 126.54 ;
   RECT 0.0 126.54 179.36 128.25 ;
   RECT 0.0 128.25 179.36 129.96 ;
   RECT 0.0 129.96 179.36 131.67 ;
   RECT 0.0 131.67 179.36 133.38 ;
   RECT 0.0 133.38 179.36 135.09 ;
   RECT 0.0 135.09 179.36 136.8 ;
   RECT 0.0 136.8 179.36 138.51 ;
   RECT 0.0 138.51 179.36 140.22 ;
   RECT 0.0 140.22 179.36 141.93 ;
   RECT 0.0 141.93 179.36 143.64 ;
   RECT 0.0 143.64 179.36 145.35 ;
   RECT 0.0 145.35 179.36 147.06 ;
   RECT 0.0 147.06 179.36 148.77 ;
   RECT 0.0 148.77 179.36 150.48 ;
   RECT 0.0 150.48 179.36 152.19 ;
   RECT 0.0 152.19 179.36 153.9 ;
   RECT 0.0 153.9 179.36 155.61 ;
   RECT 0.0 155.61 179.36 157.32 ;
   RECT 0.0 157.32 179.36 159.03 ;
   RECT 0.0 159.03 179.36 160.74 ;
   RECT 0.0 160.74 179.36 162.45 ;
   RECT 0.0 162.45 179.36 164.16 ;
   RECT 0.0 164.16 179.36 165.87 ;
   RECT 0.0 165.87 179.36 167.58 ;
   RECT 0.0 167.58 179.36 169.29 ;
   RECT 0.0 169.29 179.36 171.0 ;
   RECT 0.0 171.0 179.36 172.71 ;
   RECT 0.0 172.71 179.36 174.42 ;
   RECT 0.0 174.42 179.36 176.13 ;
   RECT 0.0 176.13 179.36 177.84 ;
   RECT 0.0 177.84 179.36 179.55 ;
   RECT 0.0 179.55 179.36 181.26 ;
   RECT 0.0 181.26 179.36 182.97 ;
   RECT 0.0 182.97 179.36 184.68 ;
   RECT 0.0 184.68 179.36 186.39 ;
   RECT 0.0 186.39 179.36 188.1 ;
   RECT 0.0 188.1 179.36 189.81 ;
   RECT 0.0 189.81 179.36 191.52 ;
   RECT 0.0 191.52 179.36 193.23 ;
   RECT 0.0 193.23 179.36 194.94 ;
   RECT 0.0 194.94 179.36 196.65 ;
   RECT 0.0 196.65 179.36 198.36 ;
  LAYER metal3 ;
   RECT 0.0 0.0 179.36 1.71 ;
   RECT 0.0 1.71 179.36 3.42 ;
   RECT 0.0 3.42 179.36 5.13 ;
   RECT 0.0 5.13 179.36 6.84 ;
   RECT 0.0 6.84 179.36 8.55 ;
   RECT 0.0 8.55 179.36 10.26 ;
   RECT 0.0 10.26 179.36 11.97 ;
   RECT 0.0 11.97 179.36 13.68 ;
   RECT 0.0 13.68 179.36 15.39 ;
   RECT 0.0 15.39 179.36 17.1 ;
   RECT 0.0 17.1 179.36 18.81 ;
   RECT 0.0 18.81 179.36 20.52 ;
   RECT 0.0 20.52 179.36 22.23 ;
   RECT 0.0 22.23 179.36 23.94 ;
   RECT 0.0 23.94 179.36 25.65 ;
   RECT 0.0 25.65 179.36 27.36 ;
   RECT 0.0 27.36 179.36 29.07 ;
   RECT 0.0 29.07 179.36 30.78 ;
   RECT 0.0 30.78 179.36 32.49 ;
   RECT 0.0 32.49 179.36 34.2 ;
   RECT 0.0 34.2 179.36 35.91 ;
   RECT 0.0 35.91 179.36 37.62 ;
   RECT 0.0 37.62 179.36 39.33 ;
   RECT 0.0 39.33 179.36 41.04 ;
   RECT 0.0 41.04 179.36 42.75 ;
   RECT 0.0 42.75 179.36 44.46 ;
   RECT 0.0 44.46 179.36 46.17 ;
   RECT 0.0 46.17 179.36 47.88 ;
   RECT 0.0 47.88 179.36 49.59 ;
   RECT 0.0 49.59 179.36 51.3 ;
   RECT 0.0 51.3 179.36 53.01 ;
   RECT 0.0 53.01 179.36 54.72 ;
   RECT 0.0 54.72 179.36 56.43 ;
   RECT 0.0 56.43 179.36 58.14 ;
   RECT 0.0 58.14 179.36 59.85 ;
   RECT 0.0 59.85 179.36 61.56 ;
   RECT 0.0 61.56 179.36 63.27 ;
   RECT 0.0 63.27 179.36 64.98 ;
   RECT 0.0 64.98 179.36 66.69 ;
   RECT 0.0 66.69 179.36 68.4 ;
   RECT 0.0 68.4 179.36 70.11 ;
   RECT 0.0 70.11 179.36 71.82 ;
   RECT 0.0 71.82 179.36 73.53 ;
   RECT 0.0 73.53 179.36 75.24 ;
   RECT 0.0 75.24 179.36 76.95 ;
   RECT 0.0 76.95 179.36 78.66 ;
   RECT 0.0 78.66 179.36 80.37 ;
   RECT 0.0 80.37 179.36 82.08 ;
   RECT 0.0 82.08 179.36 83.79 ;
   RECT 0.0 83.79 202.54 85.5 ;
   RECT 0.0 85.5 202.54 87.21 ;
   RECT 0.0 87.21 202.54 88.92 ;
   RECT 0.0 88.92 202.54 90.63 ;
   RECT 0.0 90.63 202.54 92.34 ;
   RECT 0.0 92.34 202.54 94.05 ;
   RECT 0.0 94.05 202.54 95.76 ;
   RECT 0.0 95.76 202.54 97.47 ;
   RECT 0.0 97.47 202.54 99.18 ;
   RECT 0.0 99.18 202.54 100.89 ;
   RECT 0.0 100.89 202.54 102.6 ;
   RECT 0.0 102.6 202.54 104.31 ;
   RECT 0.0 104.31 202.54 106.02 ;
   RECT 0.0 106.02 202.54 107.73 ;
   RECT 0.0 107.73 202.54 109.44 ;
   RECT 0.0 109.44 202.54 111.15 ;
   RECT 0.0 111.15 202.54 112.86 ;
   RECT 0.0 112.86 179.36 114.57 ;
   RECT 0.0 114.57 179.36 116.28 ;
   RECT 0.0 116.28 179.36 117.99 ;
   RECT 0.0 117.99 179.36 119.7 ;
   RECT 0.0 119.7 179.36 121.41 ;
   RECT 0.0 121.41 179.36 123.12 ;
   RECT 0.0 123.12 179.36 124.83 ;
   RECT 0.0 124.83 179.36 126.54 ;
   RECT 0.0 126.54 179.36 128.25 ;
   RECT 0.0 128.25 179.36 129.96 ;
   RECT 0.0 129.96 179.36 131.67 ;
   RECT 0.0 131.67 179.36 133.38 ;
   RECT 0.0 133.38 179.36 135.09 ;
   RECT 0.0 135.09 179.36 136.8 ;
   RECT 0.0 136.8 179.36 138.51 ;
   RECT 0.0 138.51 179.36 140.22 ;
   RECT 0.0 140.22 179.36 141.93 ;
   RECT 0.0 141.93 179.36 143.64 ;
   RECT 0.0 143.64 179.36 145.35 ;
   RECT 0.0 145.35 179.36 147.06 ;
   RECT 0.0 147.06 179.36 148.77 ;
   RECT 0.0 148.77 179.36 150.48 ;
   RECT 0.0 150.48 179.36 152.19 ;
   RECT 0.0 152.19 179.36 153.9 ;
   RECT 0.0 153.9 179.36 155.61 ;
   RECT 0.0 155.61 179.36 157.32 ;
   RECT 0.0 157.32 179.36 159.03 ;
   RECT 0.0 159.03 179.36 160.74 ;
   RECT 0.0 160.74 179.36 162.45 ;
   RECT 0.0 162.45 179.36 164.16 ;
   RECT 0.0 164.16 179.36 165.87 ;
   RECT 0.0 165.87 179.36 167.58 ;
   RECT 0.0 167.58 179.36 169.29 ;
   RECT 0.0 169.29 179.36 171.0 ;
   RECT 0.0 171.0 179.36 172.71 ;
   RECT 0.0 172.71 179.36 174.42 ;
   RECT 0.0 174.42 179.36 176.13 ;
   RECT 0.0 176.13 179.36 177.84 ;
   RECT 0.0 177.84 179.36 179.55 ;
   RECT 0.0 179.55 179.36 181.26 ;
   RECT 0.0 181.26 179.36 182.97 ;
   RECT 0.0 182.97 179.36 184.68 ;
   RECT 0.0 184.68 179.36 186.39 ;
   RECT 0.0 186.39 179.36 188.1 ;
   RECT 0.0 188.1 179.36 189.81 ;
   RECT 0.0 189.81 179.36 191.52 ;
   RECT 0.0 191.52 179.36 193.23 ;
   RECT 0.0 193.23 179.36 194.94 ;
   RECT 0.0 194.94 179.36 196.65 ;
   RECT 0.0 196.65 179.36 198.36 ;
  LAYER via3 ;
   RECT 0.0 0.0 179.36 1.71 ;
   RECT 0.0 1.71 179.36 3.42 ;
   RECT 0.0 3.42 179.36 5.13 ;
   RECT 0.0 5.13 179.36 6.84 ;
   RECT 0.0 6.84 179.36 8.55 ;
   RECT 0.0 8.55 179.36 10.26 ;
   RECT 0.0 10.26 179.36 11.97 ;
   RECT 0.0 11.97 179.36 13.68 ;
   RECT 0.0 13.68 179.36 15.39 ;
   RECT 0.0 15.39 179.36 17.1 ;
   RECT 0.0 17.1 179.36 18.81 ;
   RECT 0.0 18.81 179.36 20.52 ;
   RECT 0.0 20.52 179.36 22.23 ;
   RECT 0.0 22.23 179.36 23.94 ;
   RECT 0.0 23.94 179.36 25.65 ;
   RECT 0.0 25.65 179.36 27.36 ;
   RECT 0.0 27.36 179.36 29.07 ;
   RECT 0.0 29.07 179.36 30.78 ;
   RECT 0.0 30.78 179.36 32.49 ;
   RECT 0.0 32.49 179.36 34.2 ;
   RECT 0.0 34.2 179.36 35.91 ;
   RECT 0.0 35.91 179.36 37.62 ;
   RECT 0.0 37.62 179.36 39.33 ;
   RECT 0.0 39.33 179.36 41.04 ;
   RECT 0.0 41.04 179.36 42.75 ;
   RECT 0.0 42.75 179.36 44.46 ;
   RECT 0.0 44.46 179.36 46.17 ;
   RECT 0.0 46.17 179.36 47.88 ;
   RECT 0.0 47.88 179.36 49.59 ;
   RECT 0.0 49.59 179.36 51.3 ;
   RECT 0.0 51.3 179.36 53.01 ;
   RECT 0.0 53.01 179.36 54.72 ;
   RECT 0.0 54.72 179.36 56.43 ;
   RECT 0.0 56.43 179.36 58.14 ;
   RECT 0.0 58.14 179.36 59.85 ;
   RECT 0.0 59.85 179.36 61.56 ;
   RECT 0.0 61.56 179.36 63.27 ;
   RECT 0.0 63.27 179.36 64.98 ;
   RECT 0.0 64.98 179.36 66.69 ;
   RECT 0.0 66.69 179.36 68.4 ;
   RECT 0.0 68.4 179.36 70.11 ;
   RECT 0.0 70.11 179.36 71.82 ;
   RECT 0.0 71.82 179.36 73.53 ;
   RECT 0.0 73.53 179.36 75.24 ;
   RECT 0.0 75.24 179.36 76.95 ;
   RECT 0.0 76.95 179.36 78.66 ;
   RECT 0.0 78.66 179.36 80.37 ;
   RECT 0.0 80.37 179.36 82.08 ;
   RECT 0.0 82.08 179.36 83.79 ;
   RECT 0.0 83.79 202.54 85.5 ;
   RECT 0.0 85.5 202.54 87.21 ;
   RECT 0.0 87.21 202.54 88.92 ;
   RECT 0.0 88.92 202.54 90.63 ;
   RECT 0.0 90.63 202.54 92.34 ;
   RECT 0.0 92.34 202.54 94.05 ;
   RECT 0.0 94.05 202.54 95.76 ;
   RECT 0.0 95.76 202.54 97.47 ;
   RECT 0.0 97.47 202.54 99.18 ;
   RECT 0.0 99.18 202.54 100.89 ;
   RECT 0.0 100.89 202.54 102.6 ;
   RECT 0.0 102.6 202.54 104.31 ;
   RECT 0.0 104.31 202.54 106.02 ;
   RECT 0.0 106.02 202.54 107.73 ;
   RECT 0.0 107.73 202.54 109.44 ;
   RECT 0.0 109.44 202.54 111.15 ;
   RECT 0.0 111.15 202.54 112.86 ;
   RECT 0.0 112.86 179.36 114.57 ;
   RECT 0.0 114.57 179.36 116.28 ;
   RECT 0.0 116.28 179.36 117.99 ;
   RECT 0.0 117.99 179.36 119.7 ;
   RECT 0.0 119.7 179.36 121.41 ;
   RECT 0.0 121.41 179.36 123.12 ;
   RECT 0.0 123.12 179.36 124.83 ;
   RECT 0.0 124.83 179.36 126.54 ;
   RECT 0.0 126.54 179.36 128.25 ;
   RECT 0.0 128.25 179.36 129.96 ;
   RECT 0.0 129.96 179.36 131.67 ;
   RECT 0.0 131.67 179.36 133.38 ;
   RECT 0.0 133.38 179.36 135.09 ;
   RECT 0.0 135.09 179.36 136.8 ;
   RECT 0.0 136.8 179.36 138.51 ;
   RECT 0.0 138.51 179.36 140.22 ;
   RECT 0.0 140.22 179.36 141.93 ;
   RECT 0.0 141.93 179.36 143.64 ;
   RECT 0.0 143.64 179.36 145.35 ;
   RECT 0.0 145.35 179.36 147.06 ;
   RECT 0.0 147.06 179.36 148.77 ;
   RECT 0.0 148.77 179.36 150.48 ;
   RECT 0.0 150.48 179.36 152.19 ;
   RECT 0.0 152.19 179.36 153.9 ;
   RECT 0.0 153.9 179.36 155.61 ;
   RECT 0.0 155.61 179.36 157.32 ;
   RECT 0.0 157.32 179.36 159.03 ;
   RECT 0.0 159.03 179.36 160.74 ;
   RECT 0.0 160.74 179.36 162.45 ;
   RECT 0.0 162.45 179.36 164.16 ;
   RECT 0.0 164.16 179.36 165.87 ;
   RECT 0.0 165.87 179.36 167.58 ;
   RECT 0.0 167.58 179.36 169.29 ;
   RECT 0.0 169.29 179.36 171.0 ;
   RECT 0.0 171.0 179.36 172.71 ;
   RECT 0.0 172.71 179.36 174.42 ;
   RECT 0.0 174.42 179.36 176.13 ;
   RECT 0.0 176.13 179.36 177.84 ;
   RECT 0.0 177.84 179.36 179.55 ;
   RECT 0.0 179.55 179.36 181.26 ;
   RECT 0.0 181.26 179.36 182.97 ;
   RECT 0.0 182.97 179.36 184.68 ;
   RECT 0.0 184.68 179.36 186.39 ;
   RECT 0.0 186.39 179.36 188.1 ;
   RECT 0.0 188.1 179.36 189.81 ;
   RECT 0.0 189.81 179.36 191.52 ;
   RECT 0.0 191.52 179.36 193.23 ;
   RECT 0.0 193.23 179.36 194.94 ;
   RECT 0.0 194.94 179.36 196.65 ;
   RECT 0.0 196.65 179.36 198.36 ;
  LAYER metal4 ;
   RECT 0.0 0.0 179.36 1.71 ;
   RECT 0.0 1.71 179.36 3.42 ;
   RECT 0.0 3.42 179.36 5.13 ;
   RECT 0.0 5.13 179.36 6.84 ;
   RECT 0.0 6.84 179.36 8.55 ;
   RECT 0.0 8.55 179.36 10.26 ;
   RECT 0.0 10.26 179.36 11.97 ;
   RECT 0.0 11.97 179.36 13.68 ;
   RECT 0.0 13.68 179.36 15.39 ;
   RECT 0.0 15.39 179.36 17.1 ;
   RECT 0.0 17.1 179.36 18.81 ;
   RECT 0.0 18.81 179.36 20.52 ;
   RECT 0.0 20.52 179.36 22.23 ;
   RECT 0.0 22.23 179.36 23.94 ;
   RECT 0.0 23.94 179.36 25.65 ;
   RECT 0.0 25.65 179.36 27.36 ;
   RECT 0.0 27.36 179.36 29.07 ;
   RECT 0.0 29.07 179.36 30.78 ;
   RECT 0.0 30.78 179.36 32.49 ;
   RECT 0.0 32.49 179.36 34.2 ;
   RECT 0.0 34.2 179.36 35.91 ;
   RECT 0.0 35.91 179.36 37.62 ;
   RECT 0.0 37.62 179.36 39.33 ;
   RECT 0.0 39.33 179.36 41.04 ;
   RECT 0.0 41.04 179.36 42.75 ;
   RECT 0.0 42.75 179.36 44.46 ;
   RECT 0.0 44.46 179.36 46.17 ;
   RECT 0.0 46.17 179.36 47.88 ;
   RECT 0.0 47.88 179.36 49.59 ;
   RECT 0.0 49.59 179.36 51.3 ;
   RECT 0.0 51.3 179.36 53.01 ;
   RECT 0.0 53.01 179.36 54.72 ;
   RECT 0.0 54.72 179.36 56.43 ;
   RECT 0.0 56.43 179.36 58.14 ;
   RECT 0.0 58.14 179.36 59.85 ;
   RECT 0.0 59.85 179.36 61.56 ;
   RECT 0.0 61.56 179.36 63.27 ;
   RECT 0.0 63.27 179.36 64.98 ;
   RECT 0.0 64.98 179.36 66.69 ;
   RECT 0.0 66.69 179.36 68.4 ;
   RECT 0.0 68.4 179.36 70.11 ;
   RECT 0.0 70.11 179.36 71.82 ;
   RECT 0.0 71.82 179.36 73.53 ;
   RECT 0.0 73.53 179.36 75.24 ;
   RECT 0.0 75.24 179.36 76.95 ;
   RECT 0.0 76.95 179.36 78.66 ;
   RECT 0.0 78.66 179.36 80.37 ;
   RECT 0.0 80.37 179.36 82.08 ;
   RECT 0.0 82.08 179.36 83.79 ;
   RECT 0.0 83.79 202.54 85.5 ;
   RECT 0.0 85.5 202.54 87.21 ;
   RECT 0.0 87.21 202.54 88.92 ;
   RECT 0.0 88.92 202.54 90.63 ;
   RECT 0.0 90.63 202.54 92.34 ;
   RECT 0.0 92.34 202.54 94.05 ;
   RECT 0.0 94.05 202.54 95.76 ;
   RECT 0.0 95.76 202.54 97.47 ;
   RECT 0.0 97.47 202.54 99.18 ;
   RECT 0.0 99.18 202.54 100.89 ;
   RECT 0.0 100.89 202.54 102.6 ;
   RECT 0.0 102.6 202.54 104.31 ;
   RECT 0.0 104.31 202.54 106.02 ;
   RECT 0.0 106.02 202.54 107.73 ;
   RECT 0.0 107.73 202.54 109.44 ;
   RECT 0.0 109.44 202.54 111.15 ;
   RECT 0.0 111.15 202.54 112.86 ;
   RECT 0.0 112.86 179.36 114.57 ;
   RECT 0.0 114.57 179.36 116.28 ;
   RECT 0.0 116.28 179.36 117.99 ;
   RECT 0.0 117.99 179.36 119.7 ;
   RECT 0.0 119.7 179.36 121.41 ;
   RECT 0.0 121.41 179.36 123.12 ;
   RECT 0.0 123.12 179.36 124.83 ;
   RECT 0.0 124.83 179.36 126.54 ;
   RECT 0.0 126.54 179.36 128.25 ;
   RECT 0.0 128.25 179.36 129.96 ;
   RECT 0.0 129.96 179.36 131.67 ;
   RECT 0.0 131.67 179.36 133.38 ;
   RECT 0.0 133.38 179.36 135.09 ;
   RECT 0.0 135.09 179.36 136.8 ;
   RECT 0.0 136.8 179.36 138.51 ;
   RECT 0.0 138.51 179.36 140.22 ;
   RECT 0.0 140.22 179.36 141.93 ;
   RECT 0.0 141.93 179.36 143.64 ;
   RECT 0.0 143.64 179.36 145.35 ;
   RECT 0.0 145.35 179.36 147.06 ;
   RECT 0.0 147.06 179.36 148.77 ;
   RECT 0.0 148.77 179.36 150.48 ;
   RECT 0.0 150.48 179.36 152.19 ;
   RECT 0.0 152.19 179.36 153.9 ;
   RECT 0.0 153.9 179.36 155.61 ;
   RECT 0.0 155.61 179.36 157.32 ;
   RECT 0.0 157.32 179.36 159.03 ;
   RECT 0.0 159.03 179.36 160.74 ;
   RECT 0.0 160.74 179.36 162.45 ;
   RECT 0.0 162.45 179.36 164.16 ;
   RECT 0.0 164.16 179.36 165.87 ;
   RECT 0.0 165.87 179.36 167.58 ;
   RECT 0.0 167.58 179.36 169.29 ;
   RECT 0.0 169.29 179.36 171.0 ;
   RECT 0.0 171.0 179.36 172.71 ;
   RECT 0.0 172.71 179.36 174.42 ;
   RECT 0.0 174.42 179.36 176.13 ;
   RECT 0.0 176.13 179.36 177.84 ;
   RECT 0.0 177.84 179.36 179.55 ;
   RECT 0.0 179.55 179.36 181.26 ;
   RECT 0.0 181.26 179.36 182.97 ;
   RECT 0.0 182.97 179.36 184.68 ;
   RECT 0.0 184.68 179.36 186.39 ;
   RECT 0.0 186.39 179.36 188.1 ;
   RECT 0.0 188.1 179.36 189.81 ;
   RECT 0.0 189.81 179.36 191.52 ;
   RECT 0.0 191.52 179.36 193.23 ;
   RECT 0.0 193.23 179.36 194.94 ;
   RECT 0.0 194.94 179.36 196.65 ;
   RECT 0.0 196.65 179.36 198.36 ;
 END
END block_533x1044_173

MACRO block_341x369_70
 CLASS BLOCK ;
 FOREIGN block_341x369_70 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 129.58 BY 70.11 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 20.235 126.445 20.805 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 26.695 126.445 27.265 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 6.935 3.325 7.505 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 9.215 3.325 9.785 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 10.735 3.325 11.305 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 13.015 3.325 13.585 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 13.395 4.085 13.965 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 13.775 3.325 14.345 ;
  END
 END o7
 PIN o8
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 15.295 3.325 15.865 ;
  END
 END o8
 PIN o9
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 12.635 4.085 13.205 ;
  END
 END o9
 PIN o10
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 19.855 3.325 20.425 ;
  END
 END o10
 PIN o11
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 20.615 3.325 21.185 ;
  END
 END o11
 PIN o12
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 21.375 3.325 21.945 ;
  END
 END o12
 PIN o13
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 18.335 3.325 18.905 ;
  END
 END o13
 PIN o14
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 25.935 3.325 26.505 ;
  END
 END o14
 PIN o15
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 26.695 3.325 27.265 ;
  END
 END o15
 PIN o16
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 27.455 3.325 28.025 ;
  END
 END o16
 PIN o17
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 25.175 3.325 25.745 ;
  END
 END o17
 PIN o18
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 32.015 3.325 32.585 ;
  END
 END o18
 PIN o19
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 33.535 3.325 34.105 ;
  END
 END o19
 PIN o20
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 34.295 3.325 34.865 ;
  END
 END o20
 PIN o21
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 31.255 3.325 31.825 ;
  END
 END o21
 PIN o22
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 38.095 126.445 38.665 ;
  END
 END o22
 PIN o23
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 38.855 126.445 39.425 ;
  END
 END o23
 PIN o24
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 39.615 126.445 40.185 ;
  END
 END o24
 PIN o25
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 42.655 126.445 43.225 ;
  END
 END o25
 PIN o26
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 21.755 126.445 22.325 ;
  END
 END o26
 PIN o27
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 31.255 126.445 31.825 ;
  END
 END o27
 PIN o28
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 32.015 126.445 32.585 ;
  END
 END o28
 PIN o29
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 33.535 126.445 34.105 ;
  END
 END o29
 PIN o30
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 34.295 126.445 34.865 ;
  END
 END o30
 PIN o31
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 30.495 126.445 31.065 ;
  END
 END o31
 PIN o32
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 28.975 126.445 29.545 ;
  END
 END o32
 PIN o33
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 41.135 3.325 41.705 ;
  END
 END o33
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 35.815 126.445 36.385 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 43.035 125.685 43.605 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 32.395 125.685 32.965 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 35.435 125.685 36.005 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 36.955 126.445 37.525 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 36.575 125.685 37.145 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 33.915 125.685 34.485 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 30.115 125.685 30.685 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 40.375 3.325 40.945 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 8.455 3.325 9.025 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 25.935 126.445 26.505 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 25.175 126.445 25.745 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 24.415 126.445 24.985 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 34.675 125.685 35.245 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 30.875 125.685 31.445 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 40.755 126.445 41.325 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 27.455 126.445 28.025 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 38.475 125.685 39.045 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 39.995 125.685 40.565 ;
  END
 END i18
 PIN i19
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 39.235 125.685 39.805 ;
  END
 END i19
 PIN i20
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 124.355 40.375 124.925 40.945 ;
  END
 END i20
 PIN i21
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 8.455 126.445 9.025 ;
  END
 END i21
 PIN i22
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 9.215 126.445 9.785 ;
  END
 END i22
 PIN i23
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 10.735 126.445 11.305 ;
  END
 END i23
 PIN i24
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 11.495 126.445 12.065 ;
  END
 END i24
 PIN i25
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 12.255 126.445 12.825 ;
  END
 END i25
 PIN i26
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 13.015 126.445 13.585 ;
  END
 END i26
 PIN i27
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 8.075 125.685 8.645 ;
  END
 END i27
 PIN i28
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 7.695 126.445 8.265 ;
  END
 END i28
 PIN i29
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 7.315 125.685 7.885 ;
  END
 END i29
 PIN i30
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 6.935 126.445 7.505 ;
  END
 END i30
 PIN i31
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 6.555 125.685 7.125 ;
  END
 END i31
 PIN i32
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 13.775 126.445 14.345 ;
  END
 END i32
 PIN i33
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 15.295 126.445 15.865 ;
  END
 END i33
 PIN i34
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 16.055 126.445 16.625 ;
  END
 END i34
 PIN i35
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 16.815 126.445 17.385 ;
  END
 END i35
 OBS
  LAYER metal1 ;
   RECT 0 0 129.58 70.11 ;
  LAYER via1 ;
   RECT 0 0 129.58 70.11 ;
  LAYER metal2 ;
   RECT 0 0 129.58 70.11 ;
  LAYER via2 ;
   RECT 0 0 129.58 70.11 ;
  LAYER metal3 ;
   RECT 0 0 129.58 70.11 ;
  LAYER via3 ;
   RECT 0 0 129.58 70.11 ;
  LAYER metal4 ;
   RECT 0 0 129.58 70.11 ;
 END
END block_341x369_70

MACRO block_779x2502_158
 CLASS BLOCK ;
 FOREIGN block_779x2502_158 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 296.02 BY 475.38 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 465.405 269.325 465.975 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 449.065 269.325 449.635 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 283.765 269.325 284.335 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 267.425 269.325 267.995 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 251.085 269.325 251.655 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 206.625 269.325 207.195 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 190.285 269.325 190.855 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 173.945 269.325 174.515 ;
  END
 END o7
 PIN o8
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 157.605 269.325 158.175 ;
  END
 END o8
 PIN o9
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 141.265 269.325 141.835 ;
  END
 END o9
 PIN o10
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 124.925 269.325 125.495 ;
  END
 END o10
 PIN o11
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 90.345 269.325 90.915 ;
  END
 END o11
 PIN o12
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 432.725 269.325 433.295 ;
  END
 END o12
 PIN o13
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 74.005 269.325 74.575 ;
  END
 END o13
 PIN o14
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 57.665 269.325 58.235 ;
  END
 END o14
 PIN o15
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 41.325 269.325 41.895 ;
  END
 END o15
 PIN o16
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 24.985 269.325 25.555 ;
  END
 END o16
 PIN o17
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 8.645 269.325 9.215 ;
  END
 END o17
 PIN o18
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 416.385 269.325 416.955 ;
  END
 END o18
 PIN o19
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 400.045 269.325 400.615 ;
  END
 END o19
 PIN o20
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 383.705 269.325 384.275 ;
  END
 END o20
 PIN o21
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 367.365 269.325 367.935 ;
  END
 END o21
 PIN o22
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 332.785 269.325 333.355 ;
  END
 END o22
 PIN o23
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 316.445 269.325 317.015 ;
  END
 END o23
 PIN o24
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 300.105 269.325 300.675 ;
  END
 END o24
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 291.935 240.065 292.505 240.635 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 291.935 222.965 292.505 223.535 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 291.935 234.745 292.505 235.315 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 291.935 230.375 292.505 230.945 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 291.935 227.525 292.505 228.095 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 291.175 239.685 291.745 240.255 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 291.175 240.445 291.745 241.015 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 291.935 240.825 292.505 241.395 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 291.935 231.135 292.505 231.705 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 291.935 218.025 292.505 218.595 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 291.175 223.345 291.745 223.915 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 291.935 226.575 292.505 227.145 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 291.935 223.725 292.505 224.295 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 291.935 221.635 292.505 222.205 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 291.935 219.165 292.505 219.735 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 291.175 217.645 291.745 218.215 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 282.435 241.205 283.005 241.775 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 282.435 227.905 283.005 228.475 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 467.115 269.325 467.685 ;
  END
 END i18
 PIN i19
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 450.775 269.325 451.345 ;
  END
 END i19
 PIN i20
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 285.475 269.325 286.045 ;
  END
 END i20
 PIN i21
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 269.135 269.325 269.705 ;
  END
 END i21
 PIN i22
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 252.795 269.325 253.365 ;
  END
 END i22
 PIN i23
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 204.915 269.325 205.485 ;
  END
 END i23
 PIN i24
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 188.575 269.325 189.145 ;
  END
 END i24
 PIN i25
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 172.235 269.325 172.805 ;
  END
 END i25
 PIN i26
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 155.895 269.325 156.465 ;
  END
 END i26
 PIN i27
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 139.555 269.325 140.125 ;
  END
 END i27
 PIN i28
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 123.215 269.325 123.785 ;
  END
 END i28
 PIN i29
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 88.635 269.325 89.205 ;
  END
 END i29
 PIN i30
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 434.435 269.325 435.005 ;
  END
 END i30
 PIN i31
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 72.295 269.325 72.865 ;
  END
 END i31
 PIN i32
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 55.955 269.325 56.525 ;
  END
 END i32
 PIN i33
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 39.615 269.325 40.185 ;
  END
 END i33
 PIN i34
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 23.275 269.325 23.845 ;
  END
 END i34
 PIN i35
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 6.935 269.325 7.505 ;
  END
 END i35
 PIN i36
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 418.095 269.325 418.665 ;
  END
 END i36
 PIN i37
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 401.755 269.325 402.325 ;
  END
 END i37
 PIN i38
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 385.415 269.325 385.985 ;
  END
 END i38
 PIN i39
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 369.075 269.325 369.645 ;
  END
 END i39
 PIN i40
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 334.495 269.325 335.065 ;
  END
 END i40
 PIN i41
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 318.155 269.325 318.725 ;
  END
 END i41
 PIN i42
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 301.815 269.325 302.385 ;
  END
 END i42
 PIN i43
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 383.135 268.565 383.705 ;
  END
 END i43
 PIN i44
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 379.145 269.325 379.715 ;
  END
 END i44
 PIN i45
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 374.965 269.325 375.535 ;
  END
 END i45
 PIN i46
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 395.485 269.325 396.055 ;
  END
 END i46
 PIN i47
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 391.305 269.325 391.875 ;
  END
 END i47
 PIN i48
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 315.875 268.565 316.445 ;
  END
 END i48
 PIN i49
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 311.885 269.325 312.455 ;
  END
 END i49
 PIN i50
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 307.705 269.325 308.275 ;
  END
 END i50
 PIN i51
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 303.715 269.325 304.285 ;
  END
 END i51
 PIN i52
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 299.535 268.565 300.105 ;
  END
 END i52
 PIN i53
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 141.835 268.565 142.405 ;
  END
 END i53
 PIN i54
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 145.825 269.325 146.395 ;
  END
 END i54
 PIN i55
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 150.005 269.325 150.575 ;
  END
 END i55
 PIN i56
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 153.995 269.325 154.565 ;
  END
 END i56
 PIN i57
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 158.175 268.565 158.745 ;
  END
 END i57
 PIN i58
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 74.575 268.565 75.145 ;
  END
 END i58
 PIN i59
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 78.565 269.325 79.135 ;
  END
 END i59
 PIN i60
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 82.745 269.325 83.315 ;
  END
 END i60
 PIN i61
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 62.225 269.325 62.795 ;
  END
 END i61
 PIN i62
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 66.405 269.325 66.975 ;
  END
 END i62
 PIN i63
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 387.315 269.325 387.885 ;
  END
 END i63
 PIN i64
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 320.055 269.325 320.625 ;
  END
 END i64
 PIN i65
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 137.655 269.325 138.225 ;
  END
 END i65
 PIN i66
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 268.755 70.395 269.325 70.965 ;
  END
 END i66
 PIN i67
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 277.115 241.205 277.685 241.775 ;
  END
 END i67
 PIN i68
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 277.115 227.905 277.685 228.475 ;
  END
 END i68
 PIN i69
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 466.545 268.565 467.115 ;
  END
 END i69
 PIN i70
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 450.205 268.565 450.775 ;
  END
 END i70
 PIN i71
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 284.905 268.565 285.475 ;
  END
 END i71
 PIN i72
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 268.565 268.565 269.135 ;
  END
 END i72
 PIN i73
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 252.225 268.565 252.795 ;
  END
 END i73
 PIN i74
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 205.485 268.565 206.055 ;
  END
 END i74
 PIN i75
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 189.145 268.565 189.715 ;
  END
 END i75
 PIN i76
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 172.805 268.565 173.375 ;
  END
 END i76
 PIN i77
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 156.465 268.565 157.035 ;
  END
 END i77
 PIN i78
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 140.125 268.565 140.695 ;
  END
 END i78
 PIN i79
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 123.785 268.565 124.355 ;
  END
 END i79
 PIN i80
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 89.205 268.565 89.775 ;
  END
 END i80
 PIN i81
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 433.865 268.565 434.435 ;
  END
 END i81
 PIN i82
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 72.865 268.565 73.435 ;
  END
 END i82
 PIN i83
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 56.525 268.565 57.095 ;
  END
 END i83
 PIN i84
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 40.185 268.565 40.755 ;
  END
 END i84
 PIN i85
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 23.845 268.565 24.415 ;
  END
 END i85
 PIN i86
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 7.505 268.565 8.075 ;
  END
 END i86
 PIN i87
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 417.525 268.565 418.095 ;
  END
 END i87
 PIN i88
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 401.185 268.565 401.755 ;
  END
 END i88
 PIN i89
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 384.845 268.565 385.415 ;
  END
 END i89
 PIN i90
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 368.505 268.565 369.075 ;
  END
 END i90
 PIN i91
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 333.925 268.565 334.495 ;
  END
 END i91
 PIN i92
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 317.585 268.565 318.155 ;
  END
 END i92
 PIN i93
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 301.245 268.565 301.815 ;
  END
 END i93
 PIN i94
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 291.935 233.605 292.505 234.175 ;
  END
 END i94
 PIN i95
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 291.175 233.225 291.745 233.795 ;
  END
 END i95
 PIN i96
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.235 465.975 267.805 466.545 ;
  END
 END i96
 PIN i97
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.235 449.635 267.805 450.205 ;
  END
 END i97
 PIN i98
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.235 284.335 267.805 284.905 ;
  END
 END i98
 PIN i99
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.235 267.995 267.805 268.565 ;
  END
 END i99
 PIN i100
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.235 251.655 267.805 252.225 ;
  END
 END i100
 PIN i101
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.235 206.055 267.805 206.625 ;
  END
 END i101
 PIN i102
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.235 189.715 267.805 190.285 ;
  END
 END i102
 PIN i103
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.235 173.375 267.805 173.945 ;
  END
 END i103
 PIN i104
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.235 157.035 267.805 157.605 ;
  END
 END i104
 PIN i105
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.235 140.695 267.805 141.265 ;
  END
 END i105
 PIN i106
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.235 124.355 267.805 124.925 ;
  END
 END i106
 PIN i107
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.235 89.775 267.805 90.345 ;
  END
 END i107
 PIN i108
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.235 433.295 267.805 433.865 ;
  END
 END i108
 PIN i109
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.235 73.435 267.805 74.005 ;
  END
 END i109
 PIN i110
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.235 57.095 267.805 57.665 ;
  END
 END i110
 PIN i111
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.235 40.755 267.805 41.325 ;
  END
 END i111
 PIN i112
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.235 24.415 267.805 24.985 ;
  END
 END i112
 PIN i113
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.235 8.075 267.805 8.645 ;
  END
 END i113
 PIN i114
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.235 416.955 267.805 417.525 ;
  END
 END i114
 PIN i115
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.235 400.615 267.805 401.185 ;
  END
 END i115
 PIN i116
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.235 384.275 267.805 384.845 ;
  END
 END i116
 PIN i117
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.235 367.935 267.805 368.505 ;
  END
 END i117
 PIN i118
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.235 333.355 267.805 333.925 ;
  END
 END i118
 PIN i119
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.235 317.015 267.805 317.585 ;
  END
 END i119
 PIN i120
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.235 300.675 267.805 301.245 ;
  END
 END i120
 PIN i121
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 291.175 241.205 291.745 241.775 ;
  END
 END i121
 PIN i122
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 290.035 241.205 290.605 241.775 ;
  END
 END i122
 PIN i123
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 288.135 241.205 288.705 241.775 ;
  END
 END i123
 PIN i124
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 286.615 241.205 287.185 241.775 ;
  END
 END i124
 PIN i125
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 285.095 241.205 285.665 241.775 ;
  END
 END i125
 PIN i126
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 283.195 241.205 283.765 241.775 ;
  END
 END i126
 PIN i127
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 291.175 227.905 291.745 228.475 ;
  END
 END i127
 PIN i128
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 290.035 227.905 290.605 228.475 ;
  END
 END i128
 PIN i129
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 288.135 227.905 288.705 228.475 ;
  END
 END i129
 PIN i130
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 286.615 227.905 287.185 228.475 ;
  END
 END i130
 PIN i131
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 285.095 227.905 285.665 228.475 ;
  END
 END i131
 PIN i132
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 283.195 227.905 283.765 228.475 ;
  END
 END i132
 OBS
  LAYER metal1 ;
   RECT 0.0 0.0 272.84 1.71 ;
   RECT 0.0 1.71 272.84 3.42 ;
   RECT 0.0 3.42 272.84 5.13 ;
   RECT 0.0 5.13 272.84 6.84 ;
   RECT 0.0 6.84 272.84 8.55 ;
   RECT 0.0 8.55 272.84 10.26 ;
   RECT 0.0 10.26 272.84 11.97 ;
   RECT 0.0 11.97 272.84 13.68 ;
   RECT 0.0 13.68 272.84 15.39 ;
   RECT 0.0 15.39 272.84 17.1 ;
   RECT 0.0 17.1 272.84 18.81 ;
   RECT 0.0 18.81 272.84 20.52 ;
   RECT 0.0 20.52 272.84 22.23 ;
   RECT 0.0 22.23 272.84 23.94 ;
   RECT 0.0 23.94 272.84 25.65 ;
   RECT 0.0 25.65 272.84 27.36 ;
   RECT 0.0 27.36 272.84 29.07 ;
   RECT 0.0 29.07 272.84 30.78 ;
   RECT 0.0 30.78 272.84 32.49 ;
   RECT 0.0 32.49 272.84 34.2 ;
   RECT 0.0 34.2 272.84 35.91 ;
   RECT 0.0 35.91 272.84 37.62 ;
   RECT 0.0 37.62 272.84 39.33 ;
   RECT 0.0 39.33 272.84 41.04 ;
   RECT 0.0 41.04 272.84 42.75 ;
   RECT 0.0 42.75 272.84 44.46 ;
   RECT 0.0 44.46 272.84 46.17 ;
   RECT 0.0 46.17 272.84 47.88 ;
   RECT 0.0 47.88 272.84 49.59 ;
   RECT 0.0 49.59 272.84 51.3 ;
   RECT 0.0 51.3 272.84 53.01 ;
   RECT 0.0 53.01 272.84 54.72 ;
   RECT 0.0 54.72 272.84 56.43 ;
   RECT 0.0 56.43 272.84 58.14 ;
   RECT 0.0 58.14 272.84 59.85 ;
   RECT 0.0 59.85 272.84 61.56 ;
   RECT 0.0 61.56 272.84 63.27 ;
   RECT 0.0 63.27 272.84 64.98 ;
   RECT 0.0 64.98 272.84 66.69 ;
   RECT 0.0 66.69 272.84 68.4 ;
   RECT 0.0 68.4 272.84 70.11 ;
   RECT 0.0 70.11 272.84 71.82 ;
   RECT 0.0 71.82 272.84 73.53 ;
   RECT 0.0 73.53 272.84 75.24 ;
   RECT 0.0 75.24 272.84 76.95 ;
   RECT 0.0 76.95 272.84 78.66 ;
   RECT 0.0 78.66 272.84 80.37 ;
   RECT 0.0 80.37 272.84 82.08 ;
   RECT 0.0 82.08 272.84 83.79 ;
   RECT 0.0 83.79 272.84 85.5 ;
   RECT 0.0 85.5 272.84 87.21 ;
   RECT 0.0 87.21 272.84 88.92 ;
   RECT 0.0 88.92 272.84 90.63 ;
   RECT 0.0 90.63 272.84 92.34 ;
   RECT 0.0 92.34 272.84 94.05 ;
   RECT 0.0 94.05 272.84 95.76 ;
   RECT 0.0 95.76 272.84 97.47 ;
   RECT 0.0 97.47 272.84 99.18 ;
   RECT 0.0 99.18 272.84 100.89 ;
   RECT 0.0 100.89 272.84 102.6 ;
   RECT 0.0 102.6 272.84 104.31 ;
   RECT 0.0 104.31 272.84 106.02 ;
   RECT 0.0 106.02 272.84 107.73 ;
   RECT 0.0 107.73 272.84 109.44 ;
   RECT 0.0 109.44 272.84 111.15 ;
   RECT 0.0 111.15 272.84 112.86 ;
   RECT 0.0 112.86 272.84 114.57 ;
   RECT 0.0 114.57 272.84 116.28 ;
   RECT 0.0 116.28 272.84 117.99 ;
   RECT 0.0 117.99 272.84 119.7 ;
   RECT 0.0 119.7 272.84 121.41 ;
   RECT 0.0 121.41 272.84 123.12 ;
   RECT 0.0 123.12 272.84 124.83 ;
   RECT 0.0 124.83 272.84 126.54 ;
   RECT 0.0 126.54 272.84 128.25 ;
   RECT 0.0 128.25 272.84 129.96 ;
   RECT 0.0 129.96 272.84 131.67 ;
   RECT 0.0 131.67 272.84 133.38 ;
   RECT 0.0 133.38 272.84 135.09 ;
   RECT 0.0 135.09 272.84 136.8 ;
   RECT 0.0 136.8 272.84 138.51 ;
   RECT 0.0 138.51 272.84 140.22 ;
   RECT 0.0 140.22 272.84 141.93 ;
   RECT 0.0 141.93 272.84 143.64 ;
   RECT 0.0 143.64 272.84 145.35 ;
   RECT 0.0 145.35 272.84 147.06 ;
   RECT 0.0 147.06 272.84 148.77 ;
   RECT 0.0 148.77 272.84 150.48 ;
   RECT 0.0 150.48 272.84 152.19 ;
   RECT 0.0 152.19 272.84 153.9 ;
   RECT 0.0 153.9 272.84 155.61 ;
   RECT 0.0 155.61 272.84 157.32 ;
   RECT 0.0 157.32 272.84 159.03 ;
   RECT 0.0 159.03 272.84 160.74 ;
   RECT 0.0 160.74 272.84 162.45 ;
   RECT 0.0 162.45 272.84 164.16 ;
   RECT 0.0 164.16 272.84 165.87 ;
   RECT 0.0 165.87 272.84 167.58 ;
   RECT 0.0 167.58 272.84 169.29 ;
   RECT 0.0 169.29 272.84 171.0 ;
   RECT 0.0 171.0 272.84 172.71 ;
   RECT 0.0 172.71 272.84 174.42 ;
   RECT 0.0 174.42 272.84 176.13 ;
   RECT 0.0 176.13 272.84 177.84 ;
   RECT 0.0 177.84 272.84 179.55 ;
   RECT 0.0 179.55 272.84 181.26 ;
   RECT 0.0 181.26 272.84 182.97 ;
   RECT 0.0 182.97 272.84 184.68 ;
   RECT 0.0 184.68 272.84 186.39 ;
   RECT 0.0 186.39 272.84 188.1 ;
   RECT 0.0 188.1 272.84 189.81 ;
   RECT 0.0 189.81 272.84 191.52 ;
   RECT 0.0 191.52 272.84 193.23 ;
   RECT 0.0 193.23 272.84 194.94 ;
   RECT 0.0 194.94 272.84 196.65 ;
   RECT 0.0 196.65 272.84 198.36 ;
   RECT 0.0 198.36 272.84 200.07 ;
   RECT 0.0 200.07 272.84 201.78 ;
   RECT 0.0 201.78 272.84 203.49 ;
   RECT 0.0 203.49 272.84 205.2 ;
   RECT 0.0 205.2 272.84 206.91 ;
   RECT 0.0 206.91 272.84 208.62 ;
   RECT 0.0 208.62 272.84 210.33 ;
   RECT 0.0 210.33 272.84 212.04 ;
   RECT 0.0 212.04 272.84 213.75 ;
   RECT 0.0 213.75 296.02 215.46 ;
   RECT 0.0 215.46 296.02 217.17 ;
   RECT 0.0 217.17 296.02 218.88 ;
   RECT 0.0 218.88 296.02 220.59 ;
   RECT 0.0 220.59 296.02 222.3 ;
   RECT 0.0 222.3 296.02 224.01 ;
   RECT 0.0 224.01 296.02 225.72 ;
   RECT 0.0 225.72 296.02 227.43 ;
   RECT 0.0 227.43 296.02 229.14 ;
   RECT 0.0 229.14 296.02 230.85 ;
   RECT 0.0 230.85 296.02 232.56 ;
   RECT 0.0 232.56 296.02 234.27 ;
   RECT 0.0 234.27 296.02 235.98 ;
   RECT 0.0 235.98 296.02 237.69 ;
   RECT 0.0 237.69 296.02 239.4 ;
   RECT 0.0 239.4 296.02 241.11 ;
   RECT 0.0 241.11 296.02 242.82 ;
   RECT 0.0 242.82 272.84 244.53 ;
   RECT 0.0 244.53 272.84 246.24 ;
   RECT 0.0 246.24 272.84 247.95 ;
   RECT 0.0 247.95 272.84 249.66 ;
   RECT 0.0 249.66 272.84 251.37 ;
   RECT 0.0 251.37 272.84 253.08 ;
   RECT 0.0 253.08 272.84 254.79 ;
   RECT 0.0 254.79 272.84 256.5 ;
   RECT 0.0 256.5 272.84 258.21 ;
   RECT 0.0 258.21 272.84 259.92 ;
   RECT 0.0 259.92 272.84 261.63 ;
   RECT 0.0 261.63 272.84 263.34 ;
   RECT 0.0 263.34 272.84 265.05 ;
   RECT 0.0 265.05 272.84 266.76 ;
   RECT 0.0 266.76 272.84 268.47 ;
   RECT 0.0 268.47 272.84 270.18 ;
   RECT 0.0 270.18 272.84 271.89 ;
   RECT 0.0 271.89 272.84 273.6 ;
   RECT 0.0 273.6 272.84 275.31 ;
   RECT 0.0 275.31 272.84 277.02 ;
   RECT 0.0 277.02 272.84 278.73 ;
   RECT 0.0 278.73 272.84 280.44 ;
   RECT 0.0 280.44 272.84 282.15 ;
   RECT 0.0 282.15 272.84 283.86 ;
   RECT 0.0 283.86 272.84 285.57 ;
   RECT 0.0 285.57 272.84 287.28 ;
   RECT 0.0 287.28 272.84 288.99 ;
   RECT 0.0 288.99 272.84 290.7 ;
   RECT 0.0 290.7 272.84 292.41 ;
   RECT 0.0 292.41 272.84 294.12 ;
   RECT 0.0 294.12 272.84 295.83 ;
   RECT 0.0 295.83 272.84 297.54 ;
   RECT 0.0 297.54 272.84 299.25 ;
   RECT 0.0 299.25 272.84 300.96 ;
   RECT 0.0 300.96 272.84 302.67 ;
   RECT 0.0 302.67 272.84 304.38 ;
   RECT 0.0 304.38 272.84 306.09 ;
   RECT 0.0 306.09 272.84 307.8 ;
   RECT 0.0 307.8 272.84 309.51 ;
   RECT 0.0 309.51 272.84 311.22 ;
   RECT 0.0 311.22 272.84 312.93 ;
   RECT 0.0 312.93 272.84 314.64 ;
   RECT 0.0 314.64 272.84 316.35 ;
   RECT 0.0 316.35 272.84 318.06 ;
   RECT 0.0 318.06 272.84 319.77 ;
   RECT 0.0 319.77 272.84 321.48 ;
   RECT 0.0 321.48 272.84 323.19 ;
   RECT 0.0 323.19 272.84 324.9 ;
   RECT 0.0 324.9 272.84 326.61 ;
   RECT 0.0 326.61 272.84 328.32 ;
   RECT 0.0 328.32 272.84 330.03 ;
   RECT 0.0 330.03 272.84 331.74 ;
   RECT 0.0 331.74 272.84 333.45 ;
   RECT 0.0 333.45 272.84 335.16 ;
   RECT 0.0 335.16 272.84 336.87 ;
   RECT 0.0 336.87 272.84 338.58 ;
   RECT 0.0 338.58 272.84 340.29 ;
   RECT 0.0 340.29 272.84 342.0 ;
   RECT 0.0 342.0 272.84 343.71 ;
   RECT 0.0 343.71 272.84 345.42 ;
   RECT 0.0 345.42 272.84 347.13 ;
   RECT 0.0 347.13 272.84 348.84 ;
   RECT 0.0 348.84 272.84 350.55 ;
   RECT 0.0 350.55 272.84 352.26 ;
   RECT 0.0 352.26 272.84 353.97 ;
   RECT 0.0 353.97 272.84 355.68 ;
   RECT 0.0 355.68 272.84 357.39 ;
   RECT 0.0 357.39 272.84 359.1 ;
   RECT 0.0 359.1 272.84 360.81 ;
   RECT 0.0 360.81 272.84 362.52 ;
   RECT 0.0 362.52 272.84 364.23 ;
   RECT 0.0 364.23 272.84 365.94 ;
   RECT 0.0 365.94 272.84 367.65 ;
   RECT 0.0 367.65 272.84 369.36 ;
   RECT 0.0 369.36 272.84 371.07 ;
   RECT 0.0 371.07 272.84 372.78 ;
   RECT 0.0 372.78 272.84 374.49 ;
   RECT 0.0 374.49 272.84 376.2 ;
   RECT 0.0 376.2 272.84 377.91 ;
   RECT 0.0 377.91 272.84 379.62 ;
   RECT 0.0 379.62 272.84 381.33 ;
   RECT 0.0 381.33 272.84 383.04 ;
   RECT 0.0 383.04 272.84 384.75 ;
   RECT 0.0 384.75 272.84 386.46 ;
   RECT 0.0 386.46 272.84 388.17 ;
   RECT 0.0 388.17 272.84 389.88 ;
   RECT 0.0 389.88 272.84 391.59 ;
   RECT 0.0 391.59 272.84 393.3 ;
   RECT 0.0 393.3 272.84 395.01 ;
   RECT 0.0 395.01 272.84 396.72 ;
   RECT 0.0 396.72 272.84 398.43 ;
   RECT 0.0 398.43 272.84 400.14 ;
   RECT 0.0 400.14 272.84 401.85 ;
   RECT 0.0 401.85 272.84 403.56 ;
   RECT 0.0 403.56 272.84 405.27 ;
   RECT 0.0 405.27 272.84 406.98 ;
   RECT 0.0 406.98 272.84 408.69 ;
   RECT 0.0 408.69 272.84 410.4 ;
   RECT 0.0 410.4 272.84 412.11 ;
   RECT 0.0 412.11 272.84 413.82 ;
   RECT 0.0 413.82 272.84 415.53 ;
   RECT 0.0 415.53 272.84 417.24 ;
   RECT 0.0 417.24 272.84 418.95 ;
   RECT 0.0 418.95 272.84 420.66 ;
   RECT 0.0 420.66 272.84 422.37 ;
   RECT 0.0 422.37 272.84 424.08 ;
   RECT 0.0 424.08 272.84 425.79 ;
   RECT 0.0 425.79 272.84 427.5 ;
   RECT 0.0 427.5 272.84 429.21 ;
   RECT 0.0 429.21 272.84 430.92 ;
   RECT 0.0 430.92 272.84 432.63 ;
   RECT 0.0 432.63 272.84 434.34 ;
   RECT 0.0 434.34 272.84 436.05 ;
   RECT 0.0 436.05 272.84 437.76 ;
   RECT 0.0 437.76 272.84 439.47 ;
   RECT 0.0 439.47 272.84 441.18 ;
   RECT 0.0 441.18 272.84 442.89 ;
   RECT 0.0 442.89 272.84 444.6 ;
   RECT 0.0 444.6 272.84 446.31 ;
   RECT 0.0 446.31 272.84 448.02 ;
   RECT 0.0 448.02 272.84 449.73 ;
   RECT 0.0 449.73 272.84 451.44 ;
   RECT 0.0 451.44 272.84 453.15 ;
   RECT 0.0 453.15 272.84 454.86 ;
   RECT 0.0 454.86 272.84 456.57 ;
   RECT 0.0 456.57 272.84 458.28 ;
   RECT 0.0 458.28 272.84 459.99 ;
   RECT 0.0 459.99 272.84 461.7 ;
   RECT 0.0 461.7 272.84 463.41 ;
   RECT 0.0 463.41 272.84 465.12 ;
   RECT 0.0 465.12 272.84 466.83 ;
   RECT 0.0 466.83 272.84 468.54 ;
   RECT 0.0 468.54 272.84 470.25 ;
   RECT 0.0 470.25 272.84 471.96 ;
   RECT 0.0 471.96 272.84 473.67 ;
   RECT 0.0 473.67 272.84 475.38 ;
  LAYER via1 ;
   RECT 0.0 0.0 272.84 1.71 ;
   RECT 0.0 1.71 272.84 3.42 ;
   RECT 0.0 3.42 272.84 5.13 ;
   RECT 0.0 5.13 272.84 6.84 ;
   RECT 0.0 6.84 272.84 8.55 ;
   RECT 0.0 8.55 272.84 10.26 ;
   RECT 0.0 10.26 272.84 11.97 ;
   RECT 0.0 11.97 272.84 13.68 ;
   RECT 0.0 13.68 272.84 15.39 ;
   RECT 0.0 15.39 272.84 17.1 ;
   RECT 0.0 17.1 272.84 18.81 ;
   RECT 0.0 18.81 272.84 20.52 ;
   RECT 0.0 20.52 272.84 22.23 ;
   RECT 0.0 22.23 272.84 23.94 ;
   RECT 0.0 23.94 272.84 25.65 ;
   RECT 0.0 25.65 272.84 27.36 ;
   RECT 0.0 27.36 272.84 29.07 ;
   RECT 0.0 29.07 272.84 30.78 ;
   RECT 0.0 30.78 272.84 32.49 ;
   RECT 0.0 32.49 272.84 34.2 ;
   RECT 0.0 34.2 272.84 35.91 ;
   RECT 0.0 35.91 272.84 37.62 ;
   RECT 0.0 37.62 272.84 39.33 ;
   RECT 0.0 39.33 272.84 41.04 ;
   RECT 0.0 41.04 272.84 42.75 ;
   RECT 0.0 42.75 272.84 44.46 ;
   RECT 0.0 44.46 272.84 46.17 ;
   RECT 0.0 46.17 272.84 47.88 ;
   RECT 0.0 47.88 272.84 49.59 ;
   RECT 0.0 49.59 272.84 51.3 ;
   RECT 0.0 51.3 272.84 53.01 ;
   RECT 0.0 53.01 272.84 54.72 ;
   RECT 0.0 54.72 272.84 56.43 ;
   RECT 0.0 56.43 272.84 58.14 ;
   RECT 0.0 58.14 272.84 59.85 ;
   RECT 0.0 59.85 272.84 61.56 ;
   RECT 0.0 61.56 272.84 63.27 ;
   RECT 0.0 63.27 272.84 64.98 ;
   RECT 0.0 64.98 272.84 66.69 ;
   RECT 0.0 66.69 272.84 68.4 ;
   RECT 0.0 68.4 272.84 70.11 ;
   RECT 0.0 70.11 272.84 71.82 ;
   RECT 0.0 71.82 272.84 73.53 ;
   RECT 0.0 73.53 272.84 75.24 ;
   RECT 0.0 75.24 272.84 76.95 ;
   RECT 0.0 76.95 272.84 78.66 ;
   RECT 0.0 78.66 272.84 80.37 ;
   RECT 0.0 80.37 272.84 82.08 ;
   RECT 0.0 82.08 272.84 83.79 ;
   RECT 0.0 83.79 272.84 85.5 ;
   RECT 0.0 85.5 272.84 87.21 ;
   RECT 0.0 87.21 272.84 88.92 ;
   RECT 0.0 88.92 272.84 90.63 ;
   RECT 0.0 90.63 272.84 92.34 ;
   RECT 0.0 92.34 272.84 94.05 ;
   RECT 0.0 94.05 272.84 95.76 ;
   RECT 0.0 95.76 272.84 97.47 ;
   RECT 0.0 97.47 272.84 99.18 ;
   RECT 0.0 99.18 272.84 100.89 ;
   RECT 0.0 100.89 272.84 102.6 ;
   RECT 0.0 102.6 272.84 104.31 ;
   RECT 0.0 104.31 272.84 106.02 ;
   RECT 0.0 106.02 272.84 107.73 ;
   RECT 0.0 107.73 272.84 109.44 ;
   RECT 0.0 109.44 272.84 111.15 ;
   RECT 0.0 111.15 272.84 112.86 ;
   RECT 0.0 112.86 272.84 114.57 ;
   RECT 0.0 114.57 272.84 116.28 ;
   RECT 0.0 116.28 272.84 117.99 ;
   RECT 0.0 117.99 272.84 119.7 ;
   RECT 0.0 119.7 272.84 121.41 ;
   RECT 0.0 121.41 272.84 123.12 ;
   RECT 0.0 123.12 272.84 124.83 ;
   RECT 0.0 124.83 272.84 126.54 ;
   RECT 0.0 126.54 272.84 128.25 ;
   RECT 0.0 128.25 272.84 129.96 ;
   RECT 0.0 129.96 272.84 131.67 ;
   RECT 0.0 131.67 272.84 133.38 ;
   RECT 0.0 133.38 272.84 135.09 ;
   RECT 0.0 135.09 272.84 136.8 ;
   RECT 0.0 136.8 272.84 138.51 ;
   RECT 0.0 138.51 272.84 140.22 ;
   RECT 0.0 140.22 272.84 141.93 ;
   RECT 0.0 141.93 272.84 143.64 ;
   RECT 0.0 143.64 272.84 145.35 ;
   RECT 0.0 145.35 272.84 147.06 ;
   RECT 0.0 147.06 272.84 148.77 ;
   RECT 0.0 148.77 272.84 150.48 ;
   RECT 0.0 150.48 272.84 152.19 ;
   RECT 0.0 152.19 272.84 153.9 ;
   RECT 0.0 153.9 272.84 155.61 ;
   RECT 0.0 155.61 272.84 157.32 ;
   RECT 0.0 157.32 272.84 159.03 ;
   RECT 0.0 159.03 272.84 160.74 ;
   RECT 0.0 160.74 272.84 162.45 ;
   RECT 0.0 162.45 272.84 164.16 ;
   RECT 0.0 164.16 272.84 165.87 ;
   RECT 0.0 165.87 272.84 167.58 ;
   RECT 0.0 167.58 272.84 169.29 ;
   RECT 0.0 169.29 272.84 171.0 ;
   RECT 0.0 171.0 272.84 172.71 ;
   RECT 0.0 172.71 272.84 174.42 ;
   RECT 0.0 174.42 272.84 176.13 ;
   RECT 0.0 176.13 272.84 177.84 ;
   RECT 0.0 177.84 272.84 179.55 ;
   RECT 0.0 179.55 272.84 181.26 ;
   RECT 0.0 181.26 272.84 182.97 ;
   RECT 0.0 182.97 272.84 184.68 ;
   RECT 0.0 184.68 272.84 186.39 ;
   RECT 0.0 186.39 272.84 188.1 ;
   RECT 0.0 188.1 272.84 189.81 ;
   RECT 0.0 189.81 272.84 191.52 ;
   RECT 0.0 191.52 272.84 193.23 ;
   RECT 0.0 193.23 272.84 194.94 ;
   RECT 0.0 194.94 272.84 196.65 ;
   RECT 0.0 196.65 272.84 198.36 ;
   RECT 0.0 198.36 272.84 200.07 ;
   RECT 0.0 200.07 272.84 201.78 ;
   RECT 0.0 201.78 272.84 203.49 ;
   RECT 0.0 203.49 272.84 205.2 ;
   RECT 0.0 205.2 272.84 206.91 ;
   RECT 0.0 206.91 272.84 208.62 ;
   RECT 0.0 208.62 272.84 210.33 ;
   RECT 0.0 210.33 272.84 212.04 ;
   RECT 0.0 212.04 272.84 213.75 ;
   RECT 0.0 213.75 296.02 215.46 ;
   RECT 0.0 215.46 296.02 217.17 ;
   RECT 0.0 217.17 296.02 218.88 ;
   RECT 0.0 218.88 296.02 220.59 ;
   RECT 0.0 220.59 296.02 222.3 ;
   RECT 0.0 222.3 296.02 224.01 ;
   RECT 0.0 224.01 296.02 225.72 ;
   RECT 0.0 225.72 296.02 227.43 ;
   RECT 0.0 227.43 296.02 229.14 ;
   RECT 0.0 229.14 296.02 230.85 ;
   RECT 0.0 230.85 296.02 232.56 ;
   RECT 0.0 232.56 296.02 234.27 ;
   RECT 0.0 234.27 296.02 235.98 ;
   RECT 0.0 235.98 296.02 237.69 ;
   RECT 0.0 237.69 296.02 239.4 ;
   RECT 0.0 239.4 296.02 241.11 ;
   RECT 0.0 241.11 296.02 242.82 ;
   RECT 0.0 242.82 272.84 244.53 ;
   RECT 0.0 244.53 272.84 246.24 ;
   RECT 0.0 246.24 272.84 247.95 ;
   RECT 0.0 247.95 272.84 249.66 ;
   RECT 0.0 249.66 272.84 251.37 ;
   RECT 0.0 251.37 272.84 253.08 ;
   RECT 0.0 253.08 272.84 254.79 ;
   RECT 0.0 254.79 272.84 256.5 ;
   RECT 0.0 256.5 272.84 258.21 ;
   RECT 0.0 258.21 272.84 259.92 ;
   RECT 0.0 259.92 272.84 261.63 ;
   RECT 0.0 261.63 272.84 263.34 ;
   RECT 0.0 263.34 272.84 265.05 ;
   RECT 0.0 265.05 272.84 266.76 ;
   RECT 0.0 266.76 272.84 268.47 ;
   RECT 0.0 268.47 272.84 270.18 ;
   RECT 0.0 270.18 272.84 271.89 ;
   RECT 0.0 271.89 272.84 273.6 ;
   RECT 0.0 273.6 272.84 275.31 ;
   RECT 0.0 275.31 272.84 277.02 ;
   RECT 0.0 277.02 272.84 278.73 ;
   RECT 0.0 278.73 272.84 280.44 ;
   RECT 0.0 280.44 272.84 282.15 ;
   RECT 0.0 282.15 272.84 283.86 ;
   RECT 0.0 283.86 272.84 285.57 ;
   RECT 0.0 285.57 272.84 287.28 ;
   RECT 0.0 287.28 272.84 288.99 ;
   RECT 0.0 288.99 272.84 290.7 ;
   RECT 0.0 290.7 272.84 292.41 ;
   RECT 0.0 292.41 272.84 294.12 ;
   RECT 0.0 294.12 272.84 295.83 ;
   RECT 0.0 295.83 272.84 297.54 ;
   RECT 0.0 297.54 272.84 299.25 ;
   RECT 0.0 299.25 272.84 300.96 ;
   RECT 0.0 300.96 272.84 302.67 ;
   RECT 0.0 302.67 272.84 304.38 ;
   RECT 0.0 304.38 272.84 306.09 ;
   RECT 0.0 306.09 272.84 307.8 ;
   RECT 0.0 307.8 272.84 309.51 ;
   RECT 0.0 309.51 272.84 311.22 ;
   RECT 0.0 311.22 272.84 312.93 ;
   RECT 0.0 312.93 272.84 314.64 ;
   RECT 0.0 314.64 272.84 316.35 ;
   RECT 0.0 316.35 272.84 318.06 ;
   RECT 0.0 318.06 272.84 319.77 ;
   RECT 0.0 319.77 272.84 321.48 ;
   RECT 0.0 321.48 272.84 323.19 ;
   RECT 0.0 323.19 272.84 324.9 ;
   RECT 0.0 324.9 272.84 326.61 ;
   RECT 0.0 326.61 272.84 328.32 ;
   RECT 0.0 328.32 272.84 330.03 ;
   RECT 0.0 330.03 272.84 331.74 ;
   RECT 0.0 331.74 272.84 333.45 ;
   RECT 0.0 333.45 272.84 335.16 ;
   RECT 0.0 335.16 272.84 336.87 ;
   RECT 0.0 336.87 272.84 338.58 ;
   RECT 0.0 338.58 272.84 340.29 ;
   RECT 0.0 340.29 272.84 342.0 ;
   RECT 0.0 342.0 272.84 343.71 ;
   RECT 0.0 343.71 272.84 345.42 ;
   RECT 0.0 345.42 272.84 347.13 ;
   RECT 0.0 347.13 272.84 348.84 ;
   RECT 0.0 348.84 272.84 350.55 ;
   RECT 0.0 350.55 272.84 352.26 ;
   RECT 0.0 352.26 272.84 353.97 ;
   RECT 0.0 353.97 272.84 355.68 ;
   RECT 0.0 355.68 272.84 357.39 ;
   RECT 0.0 357.39 272.84 359.1 ;
   RECT 0.0 359.1 272.84 360.81 ;
   RECT 0.0 360.81 272.84 362.52 ;
   RECT 0.0 362.52 272.84 364.23 ;
   RECT 0.0 364.23 272.84 365.94 ;
   RECT 0.0 365.94 272.84 367.65 ;
   RECT 0.0 367.65 272.84 369.36 ;
   RECT 0.0 369.36 272.84 371.07 ;
   RECT 0.0 371.07 272.84 372.78 ;
   RECT 0.0 372.78 272.84 374.49 ;
   RECT 0.0 374.49 272.84 376.2 ;
   RECT 0.0 376.2 272.84 377.91 ;
   RECT 0.0 377.91 272.84 379.62 ;
   RECT 0.0 379.62 272.84 381.33 ;
   RECT 0.0 381.33 272.84 383.04 ;
   RECT 0.0 383.04 272.84 384.75 ;
   RECT 0.0 384.75 272.84 386.46 ;
   RECT 0.0 386.46 272.84 388.17 ;
   RECT 0.0 388.17 272.84 389.88 ;
   RECT 0.0 389.88 272.84 391.59 ;
   RECT 0.0 391.59 272.84 393.3 ;
   RECT 0.0 393.3 272.84 395.01 ;
   RECT 0.0 395.01 272.84 396.72 ;
   RECT 0.0 396.72 272.84 398.43 ;
   RECT 0.0 398.43 272.84 400.14 ;
   RECT 0.0 400.14 272.84 401.85 ;
   RECT 0.0 401.85 272.84 403.56 ;
   RECT 0.0 403.56 272.84 405.27 ;
   RECT 0.0 405.27 272.84 406.98 ;
   RECT 0.0 406.98 272.84 408.69 ;
   RECT 0.0 408.69 272.84 410.4 ;
   RECT 0.0 410.4 272.84 412.11 ;
   RECT 0.0 412.11 272.84 413.82 ;
   RECT 0.0 413.82 272.84 415.53 ;
   RECT 0.0 415.53 272.84 417.24 ;
   RECT 0.0 417.24 272.84 418.95 ;
   RECT 0.0 418.95 272.84 420.66 ;
   RECT 0.0 420.66 272.84 422.37 ;
   RECT 0.0 422.37 272.84 424.08 ;
   RECT 0.0 424.08 272.84 425.79 ;
   RECT 0.0 425.79 272.84 427.5 ;
   RECT 0.0 427.5 272.84 429.21 ;
   RECT 0.0 429.21 272.84 430.92 ;
   RECT 0.0 430.92 272.84 432.63 ;
   RECT 0.0 432.63 272.84 434.34 ;
   RECT 0.0 434.34 272.84 436.05 ;
   RECT 0.0 436.05 272.84 437.76 ;
   RECT 0.0 437.76 272.84 439.47 ;
   RECT 0.0 439.47 272.84 441.18 ;
   RECT 0.0 441.18 272.84 442.89 ;
   RECT 0.0 442.89 272.84 444.6 ;
   RECT 0.0 444.6 272.84 446.31 ;
   RECT 0.0 446.31 272.84 448.02 ;
   RECT 0.0 448.02 272.84 449.73 ;
   RECT 0.0 449.73 272.84 451.44 ;
   RECT 0.0 451.44 272.84 453.15 ;
   RECT 0.0 453.15 272.84 454.86 ;
   RECT 0.0 454.86 272.84 456.57 ;
   RECT 0.0 456.57 272.84 458.28 ;
   RECT 0.0 458.28 272.84 459.99 ;
   RECT 0.0 459.99 272.84 461.7 ;
   RECT 0.0 461.7 272.84 463.41 ;
   RECT 0.0 463.41 272.84 465.12 ;
   RECT 0.0 465.12 272.84 466.83 ;
   RECT 0.0 466.83 272.84 468.54 ;
   RECT 0.0 468.54 272.84 470.25 ;
   RECT 0.0 470.25 272.84 471.96 ;
   RECT 0.0 471.96 272.84 473.67 ;
   RECT 0.0 473.67 272.84 475.38 ;
  LAYER metal2 ;
   RECT 0.0 0.0 272.84 1.71 ;
   RECT 0.0 1.71 272.84 3.42 ;
   RECT 0.0 3.42 272.84 5.13 ;
   RECT 0.0 5.13 272.84 6.84 ;
   RECT 0.0 6.84 272.84 8.55 ;
   RECT 0.0 8.55 272.84 10.26 ;
   RECT 0.0 10.26 272.84 11.97 ;
   RECT 0.0 11.97 272.84 13.68 ;
   RECT 0.0 13.68 272.84 15.39 ;
   RECT 0.0 15.39 272.84 17.1 ;
   RECT 0.0 17.1 272.84 18.81 ;
   RECT 0.0 18.81 272.84 20.52 ;
   RECT 0.0 20.52 272.84 22.23 ;
   RECT 0.0 22.23 272.84 23.94 ;
   RECT 0.0 23.94 272.84 25.65 ;
   RECT 0.0 25.65 272.84 27.36 ;
   RECT 0.0 27.36 272.84 29.07 ;
   RECT 0.0 29.07 272.84 30.78 ;
   RECT 0.0 30.78 272.84 32.49 ;
   RECT 0.0 32.49 272.84 34.2 ;
   RECT 0.0 34.2 272.84 35.91 ;
   RECT 0.0 35.91 272.84 37.62 ;
   RECT 0.0 37.62 272.84 39.33 ;
   RECT 0.0 39.33 272.84 41.04 ;
   RECT 0.0 41.04 272.84 42.75 ;
   RECT 0.0 42.75 272.84 44.46 ;
   RECT 0.0 44.46 272.84 46.17 ;
   RECT 0.0 46.17 272.84 47.88 ;
   RECT 0.0 47.88 272.84 49.59 ;
   RECT 0.0 49.59 272.84 51.3 ;
   RECT 0.0 51.3 272.84 53.01 ;
   RECT 0.0 53.01 272.84 54.72 ;
   RECT 0.0 54.72 272.84 56.43 ;
   RECT 0.0 56.43 272.84 58.14 ;
   RECT 0.0 58.14 272.84 59.85 ;
   RECT 0.0 59.85 272.84 61.56 ;
   RECT 0.0 61.56 272.84 63.27 ;
   RECT 0.0 63.27 272.84 64.98 ;
   RECT 0.0 64.98 272.84 66.69 ;
   RECT 0.0 66.69 272.84 68.4 ;
   RECT 0.0 68.4 272.84 70.11 ;
   RECT 0.0 70.11 272.84 71.82 ;
   RECT 0.0 71.82 272.84 73.53 ;
   RECT 0.0 73.53 272.84 75.24 ;
   RECT 0.0 75.24 272.84 76.95 ;
   RECT 0.0 76.95 272.84 78.66 ;
   RECT 0.0 78.66 272.84 80.37 ;
   RECT 0.0 80.37 272.84 82.08 ;
   RECT 0.0 82.08 272.84 83.79 ;
   RECT 0.0 83.79 272.84 85.5 ;
   RECT 0.0 85.5 272.84 87.21 ;
   RECT 0.0 87.21 272.84 88.92 ;
   RECT 0.0 88.92 272.84 90.63 ;
   RECT 0.0 90.63 272.84 92.34 ;
   RECT 0.0 92.34 272.84 94.05 ;
   RECT 0.0 94.05 272.84 95.76 ;
   RECT 0.0 95.76 272.84 97.47 ;
   RECT 0.0 97.47 272.84 99.18 ;
   RECT 0.0 99.18 272.84 100.89 ;
   RECT 0.0 100.89 272.84 102.6 ;
   RECT 0.0 102.6 272.84 104.31 ;
   RECT 0.0 104.31 272.84 106.02 ;
   RECT 0.0 106.02 272.84 107.73 ;
   RECT 0.0 107.73 272.84 109.44 ;
   RECT 0.0 109.44 272.84 111.15 ;
   RECT 0.0 111.15 272.84 112.86 ;
   RECT 0.0 112.86 272.84 114.57 ;
   RECT 0.0 114.57 272.84 116.28 ;
   RECT 0.0 116.28 272.84 117.99 ;
   RECT 0.0 117.99 272.84 119.7 ;
   RECT 0.0 119.7 272.84 121.41 ;
   RECT 0.0 121.41 272.84 123.12 ;
   RECT 0.0 123.12 272.84 124.83 ;
   RECT 0.0 124.83 272.84 126.54 ;
   RECT 0.0 126.54 272.84 128.25 ;
   RECT 0.0 128.25 272.84 129.96 ;
   RECT 0.0 129.96 272.84 131.67 ;
   RECT 0.0 131.67 272.84 133.38 ;
   RECT 0.0 133.38 272.84 135.09 ;
   RECT 0.0 135.09 272.84 136.8 ;
   RECT 0.0 136.8 272.84 138.51 ;
   RECT 0.0 138.51 272.84 140.22 ;
   RECT 0.0 140.22 272.84 141.93 ;
   RECT 0.0 141.93 272.84 143.64 ;
   RECT 0.0 143.64 272.84 145.35 ;
   RECT 0.0 145.35 272.84 147.06 ;
   RECT 0.0 147.06 272.84 148.77 ;
   RECT 0.0 148.77 272.84 150.48 ;
   RECT 0.0 150.48 272.84 152.19 ;
   RECT 0.0 152.19 272.84 153.9 ;
   RECT 0.0 153.9 272.84 155.61 ;
   RECT 0.0 155.61 272.84 157.32 ;
   RECT 0.0 157.32 272.84 159.03 ;
   RECT 0.0 159.03 272.84 160.74 ;
   RECT 0.0 160.74 272.84 162.45 ;
   RECT 0.0 162.45 272.84 164.16 ;
   RECT 0.0 164.16 272.84 165.87 ;
   RECT 0.0 165.87 272.84 167.58 ;
   RECT 0.0 167.58 272.84 169.29 ;
   RECT 0.0 169.29 272.84 171.0 ;
   RECT 0.0 171.0 272.84 172.71 ;
   RECT 0.0 172.71 272.84 174.42 ;
   RECT 0.0 174.42 272.84 176.13 ;
   RECT 0.0 176.13 272.84 177.84 ;
   RECT 0.0 177.84 272.84 179.55 ;
   RECT 0.0 179.55 272.84 181.26 ;
   RECT 0.0 181.26 272.84 182.97 ;
   RECT 0.0 182.97 272.84 184.68 ;
   RECT 0.0 184.68 272.84 186.39 ;
   RECT 0.0 186.39 272.84 188.1 ;
   RECT 0.0 188.1 272.84 189.81 ;
   RECT 0.0 189.81 272.84 191.52 ;
   RECT 0.0 191.52 272.84 193.23 ;
   RECT 0.0 193.23 272.84 194.94 ;
   RECT 0.0 194.94 272.84 196.65 ;
   RECT 0.0 196.65 272.84 198.36 ;
   RECT 0.0 198.36 272.84 200.07 ;
   RECT 0.0 200.07 272.84 201.78 ;
   RECT 0.0 201.78 272.84 203.49 ;
   RECT 0.0 203.49 272.84 205.2 ;
   RECT 0.0 205.2 272.84 206.91 ;
   RECT 0.0 206.91 272.84 208.62 ;
   RECT 0.0 208.62 272.84 210.33 ;
   RECT 0.0 210.33 272.84 212.04 ;
   RECT 0.0 212.04 272.84 213.75 ;
   RECT 0.0 213.75 296.02 215.46 ;
   RECT 0.0 215.46 296.02 217.17 ;
   RECT 0.0 217.17 296.02 218.88 ;
   RECT 0.0 218.88 296.02 220.59 ;
   RECT 0.0 220.59 296.02 222.3 ;
   RECT 0.0 222.3 296.02 224.01 ;
   RECT 0.0 224.01 296.02 225.72 ;
   RECT 0.0 225.72 296.02 227.43 ;
   RECT 0.0 227.43 296.02 229.14 ;
   RECT 0.0 229.14 296.02 230.85 ;
   RECT 0.0 230.85 296.02 232.56 ;
   RECT 0.0 232.56 296.02 234.27 ;
   RECT 0.0 234.27 296.02 235.98 ;
   RECT 0.0 235.98 296.02 237.69 ;
   RECT 0.0 237.69 296.02 239.4 ;
   RECT 0.0 239.4 296.02 241.11 ;
   RECT 0.0 241.11 296.02 242.82 ;
   RECT 0.0 242.82 272.84 244.53 ;
   RECT 0.0 244.53 272.84 246.24 ;
   RECT 0.0 246.24 272.84 247.95 ;
   RECT 0.0 247.95 272.84 249.66 ;
   RECT 0.0 249.66 272.84 251.37 ;
   RECT 0.0 251.37 272.84 253.08 ;
   RECT 0.0 253.08 272.84 254.79 ;
   RECT 0.0 254.79 272.84 256.5 ;
   RECT 0.0 256.5 272.84 258.21 ;
   RECT 0.0 258.21 272.84 259.92 ;
   RECT 0.0 259.92 272.84 261.63 ;
   RECT 0.0 261.63 272.84 263.34 ;
   RECT 0.0 263.34 272.84 265.05 ;
   RECT 0.0 265.05 272.84 266.76 ;
   RECT 0.0 266.76 272.84 268.47 ;
   RECT 0.0 268.47 272.84 270.18 ;
   RECT 0.0 270.18 272.84 271.89 ;
   RECT 0.0 271.89 272.84 273.6 ;
   RECT 0.0 273.6 272.84 275.31 ;
   RECT 0.0 275.31 272.84 277.02 ;
   RECT 0.0 277.02 272.84 278.73 ;
   RECT 0.0 278.73 272.84 280.44 ;
   RECT 0.0 280.44 272.84 282.15 ;
   RECT 0.0 282.15 272.84 283.86 ;
   RECT 0.0 283.86 272.84 285.57 ;
   RECT 0.0 285.57 272.84 287.28 ;
   RECT 0.0 287.28 272.84 288.99 ;
   RECT 0.0 288.99 272.84 290.7 ;
   RECT 0.0 290.7 272.84 292.41 ;
   RECT 0.0 292.41 272.84 294.12 ;
   RECT 0.0 294.12 272.84 295.83 ;
   RECT 0.0 295.83 272.84 297.54 ;
   RECT 0.0 297.54 272.84 299.25 ;
   RECT 0.0 299.25 272.84 300.96 ;
   RECT 0.0 300.96 272.84 302.67 ;
   RECT 0.0 302.67 272.84 304.38 ;
   RECT 0.0 304.38 272.84 306.09 ;
   RECT 0.0 306.09 272.84 307.8 ;
   RECT 0.0 307.8 272.84 309.51 ;
   RECT 0.0 309.51 272.84 311.22 ;
   RECT 0.0 311.22 272.84 312.93 ;
   RECT 0.0 312.93 272.84 314.64 ;
   RECT 0.0 314.64 272.84 316.35 ;
   RECT 0.0 316.35 272.84 318.06 ;
   RECT 0.0 318.06 272.84 319.77 ;
   RECT 0.0 319.77 272.84 321.48 ;
   RECT 0.0 321.48 272.84 323.19 ;
   RECT 0.0 323.19 272.84 324.9 ;
   RECT 0.0 324.9 272.84 326.61 ;
   RECT 0.0 326.61 272.84 328.32 ;
   RECT 0.0 328.32 272.84 330.03 ;
   RECT 0.0 330.03 272.84 331.74 ;
   RECT 0.0 331.74 272.84 333.45 ;
   RECT 0.0 333.45 272.84 335.16 ;
   RECT 0.0 335.16 272.84 336.87 ;
   RECT 0.0 336.87 272.84 338.58 ;
   RECT 0.0 338.58 272.84 340.29 ;
   RECT 0.0 340.29 272.84 342.0 ;
   RECT 0.0 342.0 272.84 343.71 ;
   RECT 0.0 343.71 272.84 345.42 ;
   RECT 0.0 345.42 272.84 347.13 ;
   RECT 0.0 347.13 272.84 348.84 ;
   RECT 0.0 348.84 272.84 350.55 ;
   RECT 0.0 350.55 272.84 352.26 ;
   RECT 0.0 352.26 272.84 353.97 ;
   RECT 0.0 353.97 272.84 355.68 ;
   RECT 0.0 355.68 272.84 357.39 ;
   RECT 0.0 357.39 272.84 359.1 ;
   RECT 0.0 359.1 272.84 360.81 ;
   RECT 0.0 360.81 272.84 362.52 ;
   RECT 0.0 362.52 272.84 364.23 ;
   RECT 0.0 364.23 272.84 365.94 ;
   RECT 0.0 365.94 272.84 367.65 ;
   RECT 0.0 367.65 272.84 369.36 ;
   RECT 0.0 369.36 272.84 371.07 ;
   RECT 0.0 371.07 272.84 372.78 ;
   RECT 0.0 372.78 272.84 374.49 ;
   RECT 0.0 374.49 272.84 376.2 ;
   RECT 0.0 376.2 272.84 377.91 ;
   RECT 0.0 377.91 272.84 379.62 ;
   RECT 0.0 379.62 272.84 381.33 ;
   RECT 0.0 381.33 272.84 383.04 ;
   RECT 0.0 383.04 272.84 384.75 ;
   RECT 0.0 384.75 272.84 386.46 ;
   RECT 0.0 386.46 272.84 388.17 ;
   RECT 0.0 388.17 272.84 389.88 ;
   RECT 0.0 389.88 272.84 391.59 ;
   RECT 0.0 391.59 272.84 393.3 ;
   RECT 0.0 393.3 272.84 395.01 ;
   RECT 0.0 395.01 272.84 396.72 ;
   RECT 0.0 396.72 272.84 398.43 ;
   RECT 0.0 398.43 272.84 400.14 ;
   RECT 0.0 400.14 272.84 401.85 ;
   RECT 0.0 401.85 272.84 403.56 ;
   RECT 0.0 403.56 272.84 405.27 ;
   RECT 0.0 405.27 272.84 406.98 ;
   RECT 0.0 406.98 272.84 408.69 ;
   RECT 0.0 408.69 272.84 410.4 ;
   RECT 0.0 410.4 272.84 412.11 ;
   RECT 0.0 412.11 272.84 413.82 ;
   RECT 0.0 413.82 272.84 415.53 ;
   RECT 0.0 415.53 272.84 417.24 ;
   RECT 0.0 417.24 272.84 418.95 ;
   RECT 0.0 418.95 272.84 420.66 ;
   RECT 0.0 420.66 272.84 422.37 ;
   RECT 0.0 422.37 272.84 424.08 ;
   RECT 0.0 424.08 272.84 425.79 ;
   RECT 0.0 425.79 272.84 427.5 ;
   RECT 0.0 427.5 272.84 429.21 ;
   RECT 0.0 429.21 272.84 430.92 ;
   RECT 0.0 430.92 272.84 432.63 ;
   RECT 0.0 432.63 272.84 434.34 ;
   RECT 0.0 434.34 272.84 436.05 ;
   RECT 0.0 436.05 272.84 437.76 ;
   RECT 0.0 437.76 272.84 439.47 ;
   RECT 0.0 439.47 272.84 441.18 ;
   RECT 0.0 441.18 272.84 442.89 ;
   RECT 0.0 442.89 272.84 444.6 ;
   RECT 0.0 444.6 272.84 446.31 ;
   RECT 0.0 446.31 272.84 448.02 ;
   RECT 0.0 448.02 272.84 449.73 ;
   RECT 0.0 449.73 272.84 451.44 ;
   RECT 0.0 451.44 272.84 453.15 ;
   RECT 0.0 453.15 272.84 454.86 ;
   RECT 0.0 454.86 272.84 456.57 ;
   RECT 0.0 456.57 272.84 458.28 ;
   RECT 0.0 458.28 272.84 459.99 ;
   RECT 0.0 459.99 272.84 461.7 ;
   RECT 0.0 461.7 272.84 463.41 ;
   RECT 0.0 463.41 272.84 465.12 ;
   RECT 0.0 465.12 272.84 466.83 ;
   RECT 0.0 466.83 272.84 468.54 ;
   RECT 0.0 468.54 272.84 470.25 ;
   RECT 0.0 470.25 272.84 471.96 ;
   RECT 0.0 471.96 272.84 473.67 ;
   RECT 0.0 473.67 272.84 475.38 ;
  LAYER via2 ;
   RECT 0.0 0.0 272.84 1.71 ;
   RECT 0.0 1.71 272.84 3.42 ;
   RECT 0.0 3.42 272.84 5.13 ;
   RECT 0.0 5.13 272.84 6.84 ;
   RECT 0.0 6.84 272.84 8.55 ;
   RECT 0.0 8.55 272.84 10.26 ;
   RECT 0.0 10.26 272.84 11.97 ;
   RECT 0.0 11.97 272.84 13.68 ;
   RECT 0.0 13.68 272.84 15.39 ;
   RECT 0.0 15.39 272.84 17.1 ;
   RECT 0.0 17.1 272.84 18.81 ;
   RECT 0.0 18.81 272.84 20.52 ;
   RECT 0.0 20.52 272.84 22.23 ;
   RECT 0.0 22.23 272.84 23.94 ;
   RECT 0.0 23.94 272.84 25.65 ;
   RECT 0.0 25.65 272.84 27.36 ;
   RECT 0.0 27.36 272.84 29.07 ;
   RECT 0.0 29.07 272.84 30.78 ;
   RECT 0.0 30.78 272.84 32.49 ;
   RECT 0.0 32.49 272.84 34.2 ;
   RECT 0.0 34.2 272.84 35.91 ;
   RECT 0.0 35.91 272.84 37.62 ;
   RECT 0.0 37.62 272.84 39.33 ;
   RECT 0.0 39.33 272.84 41.04 ;
   RECT 0.0 41.04 272.84 42.75 ;
   RECT 0.0 42.75 272.84 44.46 ;
   RECT 0.0 44.46 272.84 46.17 ;
   RECT 0.0 46.17 272.84 47.88 ;
   RECT 0.0 47.88 272.84 49.59 ;
   RECT 0.0 49.59 272.84 51.3 ;
   RECT 0.0 51.3 272.84 53.01 ;
   RECT 0.0 53.01 272.84 54.72 ;
   RECT 0.0 54.72 272.84 56.43 ;
   RECT 0.0 56.43 272.84 58.14 ;
   RECT 0.0 58.14 272.84 59.85 ;
   RECT 0.0 59.85 272.84 61.56 ;
   RECT 0.0 61.56 272.84 63.27 ;
   RECT 0.0 63.27 272.84 64.98 ;
   RECT 0.0 64.98 272.84 66.69 ;
   RECT 0.0 66.69 272.84 68.4 ;
   RECT 0.0 68.4 272.84 70.11 ;
   RECT 0.0 70.11 272.84 71.82 ;
   RECT 0.0 71.82 272.84 73.53 ;
   RECT 0.0 73.53 272.84 75.24 ;
   RECT 0.0 75.24 272.84 76.95 ;
   RECT 0.0 76.95 272.84 78.66 ;
   RECT 0.0 78.66 272.84 80.37 ;
   RECT 0.0 80.37 272.84 82.08 ;
   RECT 0.0 82.08 272.84 83.79 ;
   RECT 0.0 83.79 272.84 85.5 ;
   RECT 0.0 85.5 272.84 87.21 ;
   RECT 0.0 87.21 272.84 88.92 ;
   RECT 0.0 88.92 272.84 90.63 ;
   RECT 0.0 90.63 272.84 92.34 ;
   RECT 0.0 92.34 272.84 94.05 ;
   RECT 0.0 94.05 272.84 95.76 ;
   RECT 0.0 95.76 272.84 97.47 ;
   RECT 0.0 97.47 272.84 99.18 ;
   RECT 0.0 99.18 272.84 100.89 ;
   RECT 0.0 100.89 272.84 102.6 ;
   RECT 0.0 102.6 272.84 104.31 ;
   RECT 0.0 104.31 272.84 106.02 ;
   RECT 0.0 106.02 272.84 107.73 ;
   RECT 0.0 107.73 272.84 109.44 ;
   RECT 0.0 109.44 272.84 111.15 ;
   RECT 0.0 111.15 272.84 112.86 ;
   RECT 0.0 112.86 272.84 114.57 ;
   RECT 0.0 114.57 272.84 116.28 ;
   RECT 0.0 116.28 272.84 117.99 ;
   RECT 0.0 117.99 272.84 119.7 ;
   RECT 0.0 119.7 272.84 121.41 ;
   RECT 0.0 121.41 272.84 123.12 ;
   RECT 0.0 123.12 272.84 124.83 ;
   RECT 0.0 124.83 272.84 126.54 ;
   RECT 0.0 126.54 272.84 128.25 ;
   RECT 0.0 128.25 272.84 129.96 ;
   RECT 0.0 129.96 272.84 131.67 ;
   RECT 0.0 131.67 272.84 133.38 ;
   RECT 0.0 133.38 272.84 135.09 ;
   RECT 0.0 135.09 272.84 136.8 ;
   RECT 0.0 136.8 272.84 138.51 ;
   RECT 0.0 138.51 272.84 140.22 ;
   RECT 0.0 140.22 272.84 141.93 ;
   RECT 0.0 141.93 272.84 143.64 ;
   RECT 0.0 143.64 272.84 145.35 ;
   RECT 0.0 145.35 272.84 147.06 ;
   RECT 0.0 147.06 272.84 148.77 ;
   RECT 0.0 148.77 272.84 150.48 ;
   RECT 0.0 150.48 272.84 152.19 ;
   RECT 0.0 152.19 272.84 153.9 ;
   RECT 0.0 153.9 272.84 155.61 ;
   RECT 0.0 155.61 272.84 157.32 ;
   RECT 0.0 157.32 272.84 159.03 ;
   RECT 0.0 159.03 272.84 160.74 ;
   RECT 0.0 160.74 272.84 162.45 ;
   RECT 0.0 162.45 272.84 164.16 ;
   RECT 0.0 164.16 272.84 165.87 ;
   RECT 0.0 165.87 272.84 167.58 ;
   RECT 0.0 167.58 272.84 169.29 ;
   RECT 0.0 169.29 272.84 171.0 ;
   RECT 0.0 171.0 272.84 172.71 ;
   RECT 0.0 172.71 272.84 174.42 ;
   RECT 0.0 174.42 272.84 176.13 ;
   RECT 0.0 176.13 272.84 177.84 ;
   RECT 0.0 177.84 272.84 179.55 ;
   RECT 0.0 179.55 272.84 181.26 ;
   RECT 0.0 181.26 272.84 182.97 ;
   RECT 0.0 182.97 272.84 184.68 ;
   RECT 0.0 184.68 272.84 186.39 ;
   RECT 0.0 186.39 272.84 188.1 ;
   RECT 0.0 188.1 272.84 189.81 ;
   RECT 0.0 189.81 272.84 191.52 ;
   RECT 0.0 191.52 272.84 193.23 ;
   RECT 0.0 193.23 272.84 194.94 ;
   RECT 0.0 194.94 272.84 196.65 ;
   RECT 0.0 196.65 272.84 198.36 ;
   RECT 0.0 198.36 272.84 200.07 ;
   RECT 0.0 200.07 272.84 201.78 ;
   RECT 0.0 201.78 272.84 203.49 ;
   RECT 0.0 203.49 272.84 205.2 ;
   RECT 0.0 205.2 272.84 206.91 ;
   RECT 0.0 206.91 272.84 208.62 ;
   RECT 0.0 208.62 272.84 210.33 ;
   RECT 0.0 210.33 272.84 212.04 ;
   RECT 0.0 212.04 272.84 213.75 ;
   RECT 0.0 213.75 296.02 215.46 ;
   RECT 0.0 215.46 296.02 217.17 ;
   RECT 0.0 217.17 296.02 218.88 ;
   RECT 0.0 218.88 296.02 220.59 ;
   RECT 0.0 220.59 296.02 222.3 ;
   RECT 0.0 222.3 296.02 224.01 ;
   RECT 0.0 224.01 296.02 225.72 ;
   RECT 0.0 225.72 296.02 227.43 ;
   RECT 0.0 227.43 296.02 229.14 ;
   RECT 0.0 229.14 296.02 230.85 ;
   RECT 0.0 230.85 296.02 232.56 ;
   RECT 0.0 232.56 296.02 234.27 ;
   RECT 0.0 234.27 296.02 235.98 ;
   RECT 0.0 235.98 296.02 237.69 ;
   RECT 0.0 237.69 296.02 239.4 ;
   RECT 0.0 239.4 296.02 241.11 ;
   RECT 0.0 241.11 296.02 242.82 ;
   RECT 0.0 242.82 272.84 244.53 ;
   RECT 0.0 244.53 272.84 246.24 ;
   RECT 0.0 246.24 272.84 247.95 ;
   RECT 0.0 247.95 272.84 249.66 ;
   RECT 0.0 249.66 272.84 251.37 ;
   RECT 0.0 251.37 272.84 253.08 ;
   RECT 0.0 253.08 272.84 254.79 ;
   RECT 0.0 254.79 272.84 256.5 ;
   RECT 0.0 256.5 272.84 258.21 ;
   RECT 0.0 258.21 272.84 259.92 ;
   RECT 0.0 259.92 272.84 261.63 ;
   RECT 0.0 261.63 272.84 263.34 ;
   RECT 0.0 263.34 272.84 265.05 ;
   RECT 0.0 265.05 272.84 266.76 ;
   RECT 0.0 266.76 272.84 268.47 ;
   RECT 0.0 268.47 272.84 270.18 ;
   RECT 0.0 270.18 272.84 271.89 ;
   RECT 0.0 271.89 272.84 273.6 ;
   RECT 0.0 273.6 272.84 275.31 ;
   RECT 0.0 275.31 272.84 277.02 ;
   RECT 0.0 277.02 272.84 278.73 ;
   RECT 0.0 278.73 272.84 280.44 ;
   RECT 0.0 280.44 272.84 282.15 ;
   RECT 0.0 282.15 272.84 283.86 ;
   RECT 0.0 283.86 272.84 285.57 ;
   RECT 0.0 285.57 272.84 287.28 ;
   RECT 0.0 287.28 272.84 288.99 ;
   RECT 0.0 288.99 272.84 290.7 ;
   RECT 0.0 290.7 272.84 292.41 ;
   RECT 0.0 292.41 272.84 294.12 ;
   RECT 0.0 294.12 272.84 295.83 ;
   RECT 0.0 295.83 272.84 297.54 ;
   RECT 0.0 297.54 272.84 299.25 ;
   RECT 0.0 299.25 272.84 300.96 ;
   RECT 0.0 300.96 272.84 302.67 ;
   RECT 0.0 302.67 272.84 304.38 ;
   RECT 0.0 304.38 272.84 306.09 ;
   RECT 0.0 306.09 272.84 307.8 ;
   RECT 0.0 307.8 272.84 309.51 ;
   RECT 0.0 309.51 272.84 311.22 ;
   RECT 0.0 311.22 272.84 312.93 ;
   RECT 0.0 312.93 272.84 314.64 ;
   RECT 0.0 314.64 272.84 316.35 ;
   RECT 0.0 316.35 272.84 318.06 ;
   RECT 0.0 318.06 272.84 319.77 ;
   RECT 0.0 319.77 272.84 321.48 ;
   RECT 0.0 321.48 272.84 323.19 ;
   RECT 0.0 323.19 272.84 324.9 ;
   RECT 0.0 324.9 272.84 326.61 ;
   RECT 0.0 326.61 272.84 328.32 ;
   RECT 0.0 328.32 272.84 330.03 ;
   RECT 0.0 330.03 272.84 331.74 ;
   RECT 0.0 331.74 272.84 333.45 ;
   RECT 0.0 333.45 272.84 335.16 ;
   RECT 0.0 335.16 272.84 336.87 ;
   RECT 0.0 336.87 272.84 338.58 ;
   RECT 0.0 338.58 272.84 340.29 ;
   RECT 0.0 340.29 272.84 342.0 ;
   RECT 0.0 342.0 272.84 343.71 ;
   RECT 0.0 343.71 272.84 345.42 ;
   RECT 0.0 345.42 272.84 347.13 ;
   RECT 0.0 347.13 272.84 348.84 ;
   RECT 0.0 348.84 272.84 350.55 ;
   RECT 0.0 350.55 272.84 352.26 ;
   RECT 0.0 352.26 272.84 353.97 ;
   RECT 0.0 353.97 272.84 355.68 ;
   RECT 0.0 355.68 272.84 357.39 ;
   RECT 0.0 357.39 272.84 359.1 ;
   RECT 0.0 359.1 272.84 360.81 ;
   RECT 0.0 360.81 272.84 362.52 ;
   RECT 0.0 362.52 272.84 364.23 ;
   RECT 0.0 364.23 272.84 365.94 ;
   RECT 0.0 365.94 272.84 367.65 ;
   RECT 0.0 367.65 272.84 369.36 ;
   RECT 0.0 369.36 272.84 371.07 ;
   RECT 0.0 371.07 272.84 372.78 ;
   RECT 0.0 372.78 272.84 374.49 ;
   RECT 0.0 374.49 272.84 376.2 ;
   RECT 0.0 376.2 272.84 377.91 ;
   RECT 0.0 377.91 272.84 379.62 ;
   RECT 0.0 379.62 272.84 381.33 ;
   RECT 0.0 381.33 272.84 383.04 ;
   RECT 0.0 383.04 272.84 384.75 ;
   RECT 0.0 384.75 272.84 386.46 ;
   RECT 0.0 386.46 272.84 388.17 ;
   RECT 0.0 388.17 272.84 389.88 ;
   RECT 0.0 389.88 272.84 391.59 ;
   RECT 0.0 391.59 272.84 393.3 ;
   RECT 0.0 393.3 272.84 395.01 ;
   RECT 0.0 395.01 272.84 396.72 ;
   RECT 0.0 396.72 272.84 398.43 ;
   RECT 0.0 398.43 272.84 400.14 ;
   RECT 0.0 400.14 272.84 401.85 ;
   RECT 0.0 401.85 272.84 403.56 ;
   RECT 0.0 403.56 272.84 405.27 ;
   RECT 0.0 405.27 272.84 406.98 ;
   RECT 0.0 406.98 272.84 408.69 ;
   RECT 0.0 408.69 272.84 410.4 ;
   RECT 0.0 410.4 272.84 412.11 ;
   RECT 0.0 412.11 272.84 413.82 ;
   RECT 0.0 413.82 272.84 415.53 ;
   RECT 0.0 415.53 272.84 417.24 ;
   RECT 0.0 417.24 272.84 418.95 ;
   RECT 0.0 418.95 272.84 420.66 ;
   RECT 0.0 420.66 272.84 422.37 ;
   RECT 0.0 422.37 272.84 424.08 ;
   RECT 0.0 424.08 272.84 425.79 ;
   RECT 0.0 425.79 272.84 427.5 ;
   RECT 0.0 427.5 272.84 429.21 ;
   RECT 0.0 429.21 272.84 430.92 ;
   RECT 0.0 430.92 272.84 432.63 ;
   RECT 0.0 432.63 272.84 434.34 ;
   RECT 0.0 434.34 272.84 436.05 ;
   RECT 0.0 436.05 272.84 437.76 ;
   RECT 0.0 437.76 272.84 439.47 ;
   RECT 0.0 439.47 272.84 441.18 ;
   RECT 0.0 441.18 272.84 442.89 ;
   RECT 0.0 442.89 272.84 444.6 ;
   RECT 0.0 444.6 272.84 446.31 ;
   RECT 0.0 446.31 272.84 448.02 ;
   RECT 0.0 448.02 272.84 449.73 ;
   RECT 0.0 449.73 272.84 451.44 ;
   RECT 0.0 451.44 272.84 453.15 ;
   RECT 0.0 453.15 272.84 454.86 ;
   RECT 0.0 454.86 272.84 456.57 ;
   RECT 0.0 456.57 272.84 458.28 ;
   RECT 0.0 458.28 272.84 459.99 ;
   RECT 0.0 459.99 272.84 461.7 ;
   RECT 0.0 461.7 272.84 463.41 ;
   RECT 0.0 463.41 272.84 465.12 ;
   RECT 0.0 465.12 272.84 466.83 ;
   RECT 0.0 466.83 272.84 468.54 ;
   RECT 0.0 468.54 272.84 470.25 ;
   RECT 0.0 470.25 272.84 471.96 ;
   RECT 0.0 471.96 272.84 473.67 ;
   RECT 0.0 473.67 272.84 475.38 ;
  LAYER metal3 ;
   RECT 0.0 0.0 272.84 1.71 ;
   RECT 0.0 1.71 272.84 3.42 ;
   RECT 0.0 3.42 272.84 5.13 ;
   RECT 0.0 5.13 272.84 6.84 ;
   RECT 0.0 6.84 272.84 8.55 ;
   RECT 0.0 8.55 272.84 10.26 ;
   RECT 0.0 10.26 272.84 11.97 ;
   RECT 0.0 11.97 272.84 13.68 ;
   RECT 0.0 13.68 272.84 15.39 ;
   RECT 0.0 15.39 272.84 17.1 ;
   RECT 0.0 17.1 272.84 18.81 ;
   RECT 0.0 18.81 272.84 20.52 ;
   RECT 0.0 20.52 272.84 22.23 ;
   RECT 0.0 22.23 272.84 23.94 ;
   RECT 0.0 23.94 272.84 25.65 ;
   RECT 0.0 25.65 272.84 27.36 ;
   RECT 0.0 27.36 272.84 29.07 ;
   RECT 0.0 29.07 272.84 30.78 ;
   RECT 0.0 30.78 272.84 32.49 ;
   RECT 0.0 32.49 272.84 34.2 ;
   RECT 0.0 34.2 272.84 35.91 ;
   RECT 0.0 35.91 272.84 37.62 ;
   RECT 0.0 37.62 272.84 39.33 ;
   RECT 0.0 39.33 272.84 41.04 ;
   RECT 0.0 41.04 272.84 42.75 ;
   RECT 0.0 42.75 272.84 44.46 ;
   RECT 0.0 44.46 272.84 46.17 ;
   RECT 0.0 46.17 272.84 47.88 ;
   RECT 0.0 47.88 272.84 49.59 ;
   RECT 0.0 49.59 272.84 51.3 ;
   RECT 0.0 51.3 272.84 53.01 ;
   RECT 0.0 53.01 272.84 54.72 ;
   RECT 0.0 54.72 272.84 56.43 ;
   RECT 0.0 56.43 272.84 58.14 ;
   RECT 0.0 58.14 272.84 59.85 ;
   RECT 0.0 59.85 272.84 61.56 ;
   RECT 0.0 61.56 272.84 63.27 ;
   RECT 0.0 63.27 272.84 64.98 ;
   RECT 0.0 64.98 272.84 66.69 ;
   RECT 0.0 66.69 272.84 68.4 ;
   RECT 0.0 68.4 272.84 70.11 ;
   RECT 0.0 70.11 272.84 71.82 ;
   RECT 0.0 71.82 272.84 73.53 ;
   RECT 0.0 73.53 272.84 75.24 ;
   RECT 0.0 75.24 272.84 76.95 ;
   RECT 0.0 76.95 272.84 78.66 ;
   RECT 0.0 78.66 272.84 80.37 ;
   RECT 0.0 80.37 272.84 82.08 ;
   RECT 0.0 82.08 272.84 83.79 ;
   RECT 0.0 83.79 272.84 85.5 ;
   RECT 0.0 85.5 272.84 87.21 ;
   RECT 0.0 87.21 272.84 88.92 ;
   RECT 0.0 88.92 272.84 90.63 ;
   RECT 0.0 90.63 272.84 92.34 ;
   RECT 0.0 92.34 272.84 94.05 ;
   RECT 0.0 94.05 272.84 95.76 ;
   RECT 0.0 95.76 272.84 97.47 ;
   RECT 0.0 97.47 272.84 99.18 ;
   RECT 0.0 99.18 272.84 100.89 ;
   RECT 0.0 100.89 272.84 102.6 ;
   RECT 0.0 102.6 272.84 104.31 ;
   RECT 0.0 104.31 272.84 106.02 ;
   RECT 0.0 106.02 272.84 107.73 ;
   RECT 0.0 107.73 272.84 109.44 ;
   RECT 0.0 109.44 272.84 111.15 ;
   RECT 0.0 111.15 272.84 112.86 ;
   RECT 0.0 112.86 272.84 114.57 ;
   RECT 0.0 114.57 272.84 116.28 ;
   RECT 0.0 116.28 272.84 117.99 ;
   RECT 0.0 117.99 272.84 119.7 ;
   RECT 0.0 119.7 272.84 121.41 ;
   RECT 0.0 121.41 272.84 123.12 ;
   RECT 0.0 123.12 272.84 124.83 ;
   RECT 0.0 124.83 272.84 126.54 ;
   RECT 0.0 126.54 272.84 128.25 ;
   RECT 0.0 128.25 272.84 129.96 ;
   RECT 0.0 129.96 272.84 131.67 ;
   RECT 0.0 131.67 272.84 133.38 ;
   RECT 0.0 133.38 272.84 135.09 ;
   RECT 0.0 135.09 272.84 136.8 ;
   RECT 0.0 136.8 272.84 138.51 ;
   RECT 0.0 138.51 272.84 140.22 ;
   RECT 0.0 140.22 272.84 141.93 ;
   RECT 0.0 141.93 272.84 143.64 ;
   RECT 0.0 143.64 272.84 145.35 ;
   RECT 0.0 145.35 272.84 147.06 ;
   RECT 0.0 147.06 272.84 148.77 ;
   RECT 0.0 148.77 272.84 150.48 ;
   RECT 0.0 150.48 272.84 152.19 ;
   RECT 0.0 152.19 272.84 153.9 ;
   RECT 0.0 153.9 272.84 155.61 ;
   RECT 0.0 155.61 272.84 157.32 ;
   RECT 0.0 157.32 272.84 159.03 ;
   RECT 0.0 159.03 272.84 160.74 ;
   RECT 0.0 160.74 272.84 162.45 ;
   RECT 0.0 162.45 272.84 164.16 ;
   RECT 0.0 164.16 272.84 165.87 ;
   RECT 0.0 165.87 272.84 167.58 ;
   RECT 0.0 167.58 272.84 169.29 ;
   RECT 0.0 169.29 272.84 171.0 ;
   RECT 0.0 171.0 272.84 172.71 ;
   RECT 0.0 172.71 272.84 174.42 ;
   RECT 0.0 174.42 272.84 176.13 ;
   RECT 0.0 176.13 272.84 177.84 ;
   RECT 0.0 177.84 272.84 179.55 ;
   RECT 0.0 179.55 272.84 181.26 ;
   RECT 0.0 181.26 272.84 182.97 ;
   RECT 0.0 182.97 272.84 184.68 ;
   RECT 0.0 184.68 272.84 186.39 ;
   RECT 0.0 186.39 272.84 188.1 ;
   RECT 0.0 188.1 272.84 189.81 ;
   RECT 0.0 189.81 272.84 191.52 ;
   RECT 0.0 191.52 272.84 193.23 ;
   RECT 0.0 193.23 272.84 194.94 ;
   RECT 0.0 194.94 272.84 196.65 ;
   RECT 0.0 196.65 272.84 198.36 ;
   RECT 0.0 198.36 272.84 200.07 ;
   RECT 0.0 200.07 272.84 201.78 ;
   RECT 0.0 201.78 272.84 203.49 ;
   RECT 0.0 203.49 272.84 205.2 ;
   RECT 0.0 205.2 272.84 206.91 ;
   RECT 0.0 206.91 272.84 208.62 ;
   RECT 0.0 208.62 272.84 210.33 ;
   RECT 0.0 210.33 272.84 212.04 ;
   RECT 0.0 212.04 272.84 213.75 ;
   RECT 0.0 213.75 296.02 215.46 ;
   RECT 0.0 215.46 296.02 217.17 ;
   RECT 0.0 217.17 296.02 218.88 ;
   RECT 0.0 218.88 296.02 220.59 ;
   RECT 0.0 220.59 296.02 222.3 ;
   RECT 0.0 222.3 296.02 224.01 ;
   RECT 0.0 224.01 296.02 225.72 ;
   RECT 0.0 225.72 296.02 227.43 ;
   RECT 0.0 227.43 296.02 229.14 ;
   RECT 0.0 229.14 296.02 230.85 ;
   RECT 0.0 230.85 296.02 232.56 ;
   RECT 0.0 232.56 296.02 234.27 ;
   RECT 0.0 234.27 296.02 235.98 ;
   RECT 0.0 235.98 296.02 237.69 ;
   RECT 0.0 237.69 296.02 239.4 ;
   RECT 0.0 239.4 296.02 241.11 ;
   RECT 0.0 241.11 296.02 242.82 ;
   RECT 0.0 242.82 272.84 244.53 ;
   RECT 0.0 244.53 272.84 246.24 ;
   RECT 0.0 246.24 272.84 247.95 ;
   RECT 0.0 247.95 272.84 249.66 ;
   RECT 0.0 249.66 272.84 251.37 ;
   RECT 0.0 251.37 272.84 253.08 ;
   RECT 0.0 253.08 272.84 254.79 ;
   RECT 0.0 254.79 272.84 256.5 ;
   RECT 0.0 256.5 272.84 258.21 ;
   RECT 0.0 258.21 272.84 259.92 ;
   RECT 0.0 259.92 272.84 261.63 ;
   RECT 0.0 261.63 272.84 263.34 ;
   RECT 0.0 263.34 272.84 265.05 ;
   RECT 0.0 265.05 272.84 266.76 ;
   RECT 0.0 266.76 272.84 268.47 ;
   RECT 0.0 268.47 272.84 270.18 ;
   RECT 0.0 270.18 272.84 271.89 ;
   RECT 0.0 271.89 272.84 273.6 ;
   RECT 0.0 273.6 272.84 275.31 ;
   RECT 0.0 275.31 272.84 277.02 ;
   RECT 0.0 277.02 272.84 278.73 ;
   RECT 0.0 278.73 272.84 280.44 ;
   RECT 0.0 280.44 272.84 282.15 ;
   RECT 0.0 282.15 272.84 283.86 ;
   RECT 0.0 283.86 272.84 285.57 ;
   RECT 0.0 285.57 272.84 287.28 ;
   RECT 0.0 287.28 272.84 288.99 ;
   RECT 0.0 288.99 272.84 290.7 ;
   RECT 0.0 290.7 272.84 292.41 ;
   RECT 0.0 292.41 272.84 294.12 ;
   RECT 0.0 294.12 272.84 295.83 ;
   RECT 0.0 295.83 272.84 297.54 ;
   RECT 0.0 297.54 272.84 299.25 ;
   RECT 0.0 299.25 272.84 300.96 ;
   RECT 0.0 300.96 272.84 302.67 ;
   RECT 0.0 302.67 272.84 304.38 ;
   RECT 0.0 304.38 272.84 306.09 ;
   RECT 0.0 306.09 272.84 307.8 ;
   RECT 0.0 307.8 272.84 309.51 ;
   RECT 0.0 309.51 272.84 311.22 ;
   RECT 0.0 311.22 272.84 312.93 ;
   RECT 0.0 312.93 272.84 314.64 ;
   RECT 0.0 314.64 272.84 316.35 ;
   RECT 0.0 316.35 272.84 318.06 ;
   RECT 0.0 318.06 272.84 319.77 ;
   RECT 0.0 319.77 272.84 321.48 ;
   RECT 0.0 321.48 272.84 323.19 ;
   RECT 0.0 323.19 272.84 324.9 ;
   RECT 0.0 324.9 272.84 326.61 ;
   RECT 0.0 326.61 272.84 328.32 ;
   RECT 0.0 328.32 272.84 330.03 ;
   RECT 0.0 330.03 272.84 331.74 ;
   RECT 0.0 331.74 272.84 333.45 ;
   RECT 0.0 333.45 272.84 335.16 ;
   RECT 0.0 335.16 272.84 336.87 ;
   RECT 0.0 336.87 272.84 338.58 ;
   RECT 0.0 338.58 272.84 340.29 ;
   RECT 0.0 340.29 272.84 342.0 ;
   RECT 0.0 342.0 272.84 343.71 ;
   RECT 0.0 343.71 272.84 345.42 ;
   RECT 0.0 345.42 272.84 347.13 ;
   RECT 0.0 347.13 272.84 348.84 ;
   RECT 0.0 348.84 272.84 350.55 ;
   RECT 0.0 350.55 272.84 352.26 ;
   RECT 0.0 352.26 272.84 353.97 ;
   RECT 0.0 353.97 272.84 355.68 ;
   RECT 0.0 355.68 272.84 357.39 ;
   RECT 0.0 357.39 272.84 359.1 ;
   RECT 0.0 359.1 272.84 360.81 ;
   RECT 0.0 360.81 272.84 362.52 ;
   RECT 0.0 362.52 272.84 364.23 ;
   RECT 0.0 364.23 272.84 365.94 ;
   RECT 0.0 365.94 272.84 367.65 ;
   RECT 0.0 367.65 272.84 369.36 ;
   RECT 0.0 369.36 272.84 371.07 ;
   RECT 0.0 371.07 272.84 372.78 ;
   RECT 0.0 372.78 272.84 374.49 ;
   RECT 0.0 374.49 272.84 376.2 ;
   RECT 0.0 376.2 272.84 377.91 ;
   RECT 0.0 377.91 272.84 379.62 ;
   RECT 0.0 379.62 272.84 381.33 ;
   RECT 0.0 381.33 272.84 383.04 ;
   RECT 0.0 383.04 272.84 384.75 ;
   RECT 0.0 384.75 272.84 386.46 ;
   RECT 0.0 386.46 272.84 388.17 ;
   RECT 0.0 388.17 272.84 389.88 ;
   RECT 0.0 389.88 272.84 391.59 ;
   RECT 0.0 391.59 272.84 393.3 ;
   RECT 0.0 393.3 272.84 395.01 ;
   RECT 0.0 395.01 272.84 396.72 ;
   RECT 0.0 396.72 272.84 398.43 ;
   RECT 0.0 398.43 272.84 400.14 ;
   RECT 0.0 400.14 272.84 401.85 ;
   RECT 0.0 401.85 272.84 403.56 ;
   RECT 0.0 403.56 272.84 405.27 ;
   RECT 0.0 405.27 272.84 406.98 ;
   RECT 0.0 406.98 272.84 408.69 ;
   RECT 0.0 408.69 272.84 410.4 ;
   RECT 0.0 410.4 272.84 412.11 ;
   RECT 0.0 412.11 272.84 413.82 ;
   RECT 0.0 413.82 272.84 415.53 ;
   RECT 0.0 415.53 272.84 417.24 ;
   RECT 0.0 417.24 272.84 418.95 ;
   RECT 0.0 418.95 272.84 420.66 ;
   RECT 0.0 420.66 272.84 422.37 ;
   RECT 0.0 422.37 272.84 424.08 ;
   RECT 0.0 424.08 272.84 425.79 ;
   RECT 0.0 425.79 272.84 427.5 ;
   RECT 0.0 427.5 272.84 429.21 ;
   RECT 0.0 429.21 272.84 430.92 ;
   RECT 0.0 430.92 272.84 432.63 ;
   RECT 0.0 432.63 272.84 434.34 ;
   RECT 0.0 434.34 272.84 436.05 ;
   RECT 0.0 436.05 272.84 437.76 ;
   RECT 0.0 437.76 272.84 439.47 ;
   RECT 0.0 439.47 272.84 441.18 ;
   RECT 0.0 441.18 272.84 442.89 ;
   RECT 0.0 442.89 272.84 444.6 ;
   RECT 0.0 444.6 272.84 446.31 ;
   RECT 0.0 446.31 272.84 448.02 ;
   RECT 0.0 448.02 272.84 449.73 ;
   RECT 0.0 449.73 272.84 451.44 ;
   RECT 0.0 451.44 272.84 453.15 ;
   RECT 0.0 453.15 272.84 454.86 ;
   RECT 0.0 454.86 272.84 456.57 ;
   RECT 0.0 456.57 272.84 458.28 ;
   RECT 0.0 458.28 272.84 459.99 ;
   RECT 0.0 459.99 272.84 461.7 ;
   RECT 0.0 461.7 272.84 463.41 ;
   RECT 0.0 463.41 272.84 465.12 ;
   RECT 0.0 465.12 272.84 466.83 ;
   RECT 0.0 466.83 272.84 468.54 ;
   RECT 0.0 468.54 272.84 470.25 ;
   RECT 0.0 470.25 272.84 471.96 ;
   RECT 0.0 471.96 272.84 473.67 ;
   RECT 0.0 473.67 272.84 475.38 ;
  LAYER via3 ;
   RECT 0.0 0.0 272.84 1.71 ;
   RECT 0.0 1.71 272.84 3.42 ;
   RECT 0.0 3.42 272.84 5.13 ;
   RECT 0.0 5.13 272.84 6.84 ;
   RECT 0.0 6.84 272.84 8.55 ;
   RECT 0.0 8.55 272.84 10.26 ;
   RECT 0.0 10.26 272.84 11.97 ;
   RECT 0.0 11.97 272.84 13.68 ;
   RECT 0.0 13.68 272.84 15.39 ;
   RECT 0.0 15.39 272.84 17.1 ;
   RECT 0.0 17.1 272.84 18.81 ;
   RECT 0.0 18.81 272.84 20.52 ;
   RECT 0.0 20.52 272.84 22.23 ;
   RECT 0.0 22.23 272.84 23.94 ;
   RECT 0.0 23.94 272.84 25.65 ;
   RECT 0.0 25.65 272.84 27.36 ;
   RECT 0.0 27.36 272.84 29.07 ;
   RECT 0.0 29.07 272.84 30.78 ;
   RECT 0.0 30.78 272.84 32.49 ;
   RECT 0.0 32.49 272.84 34.2 ;
   RECT 0.0 34.2 272.84 35.91 ;
   RECT 0.0 35.91 272.84 37.62 ;
   RECT 0.0 37.62 272.84 39.33 ;
   RECT 0.0 39.33 272.84 41.04 ;
   RECT 0.0 41.04 272.84 42.75 ;
   RECT 0.0 42.75 272.84 44.46 ;
   RECT 0.0 44.46 272.84 46.17 ;
   RECT 0.0 46.17 272.84 47.88 ;
   RECT 0.0 47.88 272.84 49.59 ;
   RECT 0.0 49.59 272.84 51.3 ;
   RECT 0.0 51.3 272.84 53.01 ;
   RECT 0.0 53.01 272.84 54.72 ;
   RECT 0.0 54.72 272.84 56.43 ;
   RECT 0.0 56.43 272.84 58.14 ;
   RECT 0.0 58.14 272.84 59.85 ;
   RECT 0.0 59.85 272.84 61.56 ;
   RECT 0.0 61.56 272.84 63.27 ;
   RECT 0.0 63.27 272.84 64.98 ;
   RECT 0.0 64.98 272.84 66.69 ;
   RECT 0.0 66.69 272.84 68.4 ;
   RECT 0.0 68.4 272.84 70.11 ;
   RECT 0.0 70.11 272.84 71.82 ;
   RECT 0.0 71.82 272.84 73.53 ;
   RECT 0.0 73.53 272.84 75.24 ;
   RECT 0.0 75.24 272.84 76.95 ;
   RECT 0.0 76.95 272.84 78.66 ;
   RECT 0.0 78.66 272.84 80.37 ;
   RECT 0.0 80.37 272.84 82.08 ;
   RECT 0.0 82.08 272.84 83.79 ;
   RECT 0.0 83.79 272.84 85.5 ;
   RECT 0.0 85.5 272.84 87.21 ;
   RECT 0.0 87.21 272.84 88.92 ;
   RECT 0.0 88.92 272.84 90.63 ;
   RECT 0.0 90.63 272.84 92.34 ;
   RECT 0.0 92.34 272.84 94.05 ;
   RECT 0.0 94.05 272.84 95.76 ;
   RECT 0.0 95.76 272.84 97.47 ;
   RECT 0.0 97.47 272.84 99.18 ;
   RECT 0.0 99.18 272.84 100.89 ;
   RECT 0.0 100.89 272.84 102.6 ;
   RECT 0.0 102.6 272.84 104.31 ;
   RECT 0.0 104.31 272.84 106.02 ;
   RECT 0.0 106.02 272.84 107.73 ;
   RECT 0.0 107.73 272.84 109.44 ;
   RECT 0.0 109.44 272.84 111.15 ;
   RECT 0.0 111.15 272.84 112.86 ;
   RECT 0.0 112.86 272.84 114.57 ;
   RECT 0.0 114.57 272.84 116.28 ;
   RECT 0.0 116.28 272.84 117.99 ;
   RECT 0.0 117.99 272.84 119.7 ;
   RECT 0.0 119.7 272.84 121.41 ;
   RECT 0.0 121.41 272.84 123.12 ;
   RECT 0.0 123.12 272.84 124.83 ;
   RECT 0.0 124.83 272.84 126.54 ;
   RECT 0.0 126.54 272.84 128.25 ;
   RECT 0.0 128.25 272.84 129.96 ;
   RECT 0.0 129.96 272.84 131.67 ;
   RECT 0.0 131.67 272.84 133.38 ;
   RECT 0.0 133.38 272.84 135.09 ;
   RECT 0.0 135.09 272.84 136.8 ;
   RECT 0.0 136.8 272.84 138.51 ;
   RECT 0.0 138.51 272.84 140.22 ;
   RECT 0.0 140.22 272.84 141.93 ;
   RECT 0.0 141.93 272.84 143.64 ;
   RECT 0.0 143.64 272.84 145.35 ;
   RECT 0.0 145.35 272.84 147.06 ;
   RECT 0.0 147.06 272.84 148.77 ;
   RECT 0.0 148.77 272.84 150.48 ;
   RECT 0.0 150.48 272.84 152.19 ;
   RECT 0.0 152.19 272.84 153.9 ;
   RECT 0.0 153.9 272.84 155.61 ;
   RECT 0.0 155.61 272.84 157.32 ;
   RECT 0.0 157.32 272.84 159.03 ;
   RECT 0.0 159.03 272.84 160.74 ;
   RECT 0.0 160.74 272.84 162.45 ;
   RECT 0.0 162.45 272.84 164.16 ;
   RECT 0.0 164.16 272.84 165.87 ;
   RECT 0.0 165.87 272.84 167.58 ;
   RECT 0.0 167.58 272.84 169.29 ;
   RECT 0.0 169.29 272.84 171.0 ;
   RECT 0.0 171.0 272.84 172.71 ;
   RECT 0.0 172.71 272.84 174.42 ;
   RECT 0.0 174.42 272.84 176.13 ;
   RECT 0.0 176.13 272.84 177.84 ;
   RECT 0.0 177.84 272.84 179.55 ;
   RECT 0.0 179.55 272.84 181.26 ;
   RECT 0.0 181.26 272.84 182.97 ;
   RECT 0.0 182.97 272.84 184.68 ;
   RECT 0.0 184.68 272.84 186.39 ;
   RECT 0.0 186.39 272.84 188.1 ;
   RECT 0.0 188.1 272.84 189.81 ;
   RECT 0.0 189.81 272.84 191.52 ;
   RECT 0.0 191.52 272.84 193.23 ;
   RECT 0.0 193.23 272.84 194.94 ;
   RECT 0.0 194.94 272.84 196.65 ;
   RECT 0.0 196.65 272.84 198.36 ;
   RECT 0.0 198.36 272.84 200.07 ;
   RECT 0.0 200.07 272.84 201.78 ;
   RECT 0.0 201.78 272.84 203.49 ;
   RECT 0.0 203.49 272.84 205.2 ;
   RECT 0.0 205.2 272.84 206.91 ;
   RECT 0.0 206.91 272.84 208.62 ;
   RECT 0.0 208.62 272.84 210.33 ;
   RECT 0.0 210.33 272.84 212.04 ;
   RECT 0.0 212.04 272.84 213.75 ;
   RECT 0.0 213.75 296.02 215.46 ;
   RECT 0.0 215.46 296.02 217.17 ;
   RECT 0.0 217.17 296.02 218.88 ;
   RECT 0.0 218.88 296.02 220.59 ;
   RECT 0.0 220.59 296.02 222.3 ;
   RECT 0.0 222.3 296.02 224.01 ;
   RECT 0.0 224.01 296.02 225.72 ;
   RECT 0.0 225.72 296.02 227.43 ;
   RECT 0.0 227.43 296.02 229.14 ;
   RECT 0.0 229.14 296.02 230.85 ;
   RECT 0.0 230.85 296.02 232.56 ;
   RECT 0.0 232.56 296.02 234.27 ;
   RECT 0.0 234.27 296.02 235.98 ;
   RECT 0.0 235.98 296.02 237.69 ;
   RECT 0.0 237.69 296.02 239.4 ;
   RECT 0.0 239.4 296.02 241.11 ;
   RECT 0.0 241.11 296.02 242.82 ;
   RECT 0.0 242.82 272.84 244.53 ;
   RECT 0.0 244.53 272.84 246.24 ;
   RECT 0.0 246.24 272.84 247.95 ;
   RECT 0.0 247.95 272.84 249.66 ;
   RECT 0.0 249.66 272.84 251.37 ;
   RECT 0.0 251.37 272.84 253.08 ;
   RECT 0.0 253.08 272.84 254.79 ;
   RECT 0.0 254.79 272.84 256.5 ;
   RECT 0.0 256.5 272.84 258.21 ;
   RECT 0.0 258.21 272.84 259.92 ;
   RECT 0.0 259.92 272.84 261.63 ;
   RECT 0.0 261.63 272.84 263.34 ;
   RECT 0.0 263.34 272.84 265.05 ;
   RECT 0.0 265.05 272.84 266.76 ;
   RECT 0.0 266.76 272.84 268.47 ;
   RECT 0.0 268.47 272.84 270.18 ;
   RECT 0.0 270.18 272.84 271.89 ;
   RECT 0.0 271.89 272.84 273.6 ;
   RECT 0.0 273.6 272.84 275.31 ;
   RECT 0.0 275.31 272.84 277.02 ;
   RECT 0.0 277.02 272.84 278.73 ;
   RECT 0.0 278.73 272.84 280.44 ;
   RECT 0.0 280.44 272.84 282.15 ;
   RECT 0.0 282.15 272.84 283.86 ;
   RECT 0.0 283.86 272.84 285.57 ;
   RECT 0.0 285.57 272.84 287.28 ;
   RECT 0.0 287.28 272.84 288.99 ;
   RECT 0.0 288.99 272.84 290.7 ;
   RECT 0.0 290.7 272.84 292.41 ;
   RECT 0.0 292.41 272.84 294.12 ;
   RECT 0.0 294.12 272.84 295.83 ;
   RECT 0.0 295.83 272.84 297.54 ;
   RECT 0.0 297.54 272.84 299.25 ;
   RECT 0.0 299.25 272.84 300.96 ;
   RECT 0.0 300.96 272.84 302.67 ;
   RECT 0.0 302.67 272.84 304.38 ;
   RECT 0.0 304.38 272.84 306.09 ;
   RECT 0.0 306.09 272.84 307.8 ;
   RECT 0.0 307.8 272.84 309.51 ;
   RECT 0.0 309.51 272.84 311.22 ;
   RECT 0.0 311.22 272.84 312.93 ;
   RECT 0.0 312.93 272.84 314.64 ;
   RECT 0.0 314.64 272.84 316.35 ;
   RECT 0.0 316.35 272.84 318.06 ;
   RECT 0.0 318.06 272.84 319.77 ;
   RECT 0.0 319.77 272.84 321.48 ;
   RECT 0.0 321.48 272.84 323.19 ;
   RECT 0.0 323.19 272.84 324.9 ;
   RECT 0.0 324.9 272.84 326.61 ;
   RECT 0.0 326.61 272.84 328.32 ;
   RECT 0.0 328.32 272.84 330.03 ;
   RECT 0.0 330.03 272.84 331.74 ;
   RECT 0.0 331.74 272.84 333.45 ;
   RECT 0.0 333.45 272.84 335.16 ;
   RECT 0.0 335.16 272.84 336.87 ;
   RECT 0.0 336.87 272.84 338.58 ;
   RECT 0.0 338.58 272.84 340.29 ;
   RECT 0.0 340.29 272.84 342.0 ;
   RECT 0.0 342.0 272.84 343.71 ;
   RECT 0.0 343.71 272.84 345.42 ;
   RECT 0.0 345.42 272.84 347.13 ;
   RECT 0.0 347.13 272.84 348.84 ;
   RECT 0.0 348.84 272.84 350.55 ;
   RECT 0.0 350.55 272.84 352.26 ;
   RECT 0.0 352.26 272.84 353.97 ;
   RECT 0.0 353.97 272.84 355.68 ;
   RECT 0.0 355.68 272.84 357.39 ;
   RECT 0.0 357.39 272.84 359.1 ;
   RECT 0.0 359.1 272.84 360.81 ;
   RECT 0.0 360.81 272.84 362.52 ;
   RECT 0.0 362.52 272.84 364.23 ;
   RECT 0.0 364.23 272.84 365.94 ;
   RECT 0.0 365.94 272.84 367.65 ;
   RECT 0.0 367.65 272.84 369.36 ;
   RECT 0.0 369.36 272.84 371.07 ;
   RECT 0.0 371.07 272.84 372.78 ;
   RECT 0.0 372.78 272.84 374.49 ;
   RECT 0.0 374.49 272.84 376.2 ;
   RECT 0.0 376.2 272.84 377.91 ;
   RECT 0.0 377.91 272.84 379.62 ;
   RECT 0.0 379.62 272.84 381.33 ;
   RECT 0.0 381.33 272.84 383.04 ;
   RECT 0.0 383.04 272.84 384.75 ;
   RECT 0.0 384.75 272.84 386.46 ;
   RECT 0.0 386.46 272.84 388.17 ;
   RECT 0.0 388.17 272.84 389.88 ;
   RECT 0.0 389.88 272.84 391.59 ;
   RECT 0.0 391.59 272.84 393.3 ;
   RECT 0.0 393.3 272.84 395.01 ;
   RECT 0.0 395.01 272.84 396.72 ;
   RECT 0.0 396.72 272.84 398.43 ;
   RECT 0.0 398.43 272.84 400.14 ;
   RECT 0.0 400.14 272.84 401.85 ;
   RECT 0.0 401.85 272.84 403.56 ;
   RECT 0.0 403.56 272.84 405.27 ;
   RECT 0.0 405.27 272.84 406.98 ;
   RECT 0.0 406.98 272.84 408.69 ;
   RECT 0.0 408.69 272.84 410.4 ;
   RECT 0.0 410.4 272.84 412.11 ;
   RECT 0.0 412.11 272.84 413.82 ;
   RECT 0.0 413.82 272.84 415.53 ;
   RECT 0.0 415.53 272.84 417.24 ;
   RECT 0.0 417.24 272.84 418.95 ;
   RECT 0.0 418.95 272.84 420.66 ;
   RECT 0.0 420.66 272.84 422.37 ;
   RECT 0.0 422.37 272.84 424.08 ;
   RECT 0.0 424.08 272.84 425.79 ;
   RECT 0.0 425.79 272.84 427.5 ;
   RECT 0.0 427.5 272.84 429.21 ;
   RECT 0.0 429.21 272.84 430.92 ;
   RECT 0.0 430.92 272.84 432.63 ;
   RECT 0.0 432.63 272.84 434.34 ;
   RECT 0.0 434.34 272.84 436.05 ;
   RECT 0.0 436.05 272.84 437.76 ;
   RECT 0.0 437.76 272.84 439.47 ;
   RECT 0.0 439.47 272.84 441.18 ;
   RECT 0.0 441.18 272.84 442.89 ;
   RECT 0.0 442.89 272.84 444.6 ;
   RECT 0.0 444.6 272.84 446.31 ;
   RECT 0.0 446.31 272.84 448.02 ;
   RECT 0.0 448.02 272.84 449.73 ;
   RECT 0.0 449.73 272.84 451.44 ;
   RECT 0.0 451.44 272.84 453.15 ;
   RECT 0.0 453.15 272.84 454.86 ;
   RECT 0.0 454.86 272.84 456.57 ;
   RECT 0.0 456.57 272.84 458.28 ;
   RECT 0.0 458.28 272.84 459.99 ;
   RECT 0.0 459.99 272.84 461.7 ;
   RECT 0.0 461.7 272.84 463.41 ;
   RECT 0.0 463.41 272.84 465.12 ;
   RECT 0.0 465.12 272.84 466.83 ;
   RECT 0.0 466.83 272.84 468.54 ;
   RECT 0.0 468.54 272.84 470.25 ;
   RECT 0.0 470.25 272.84 471.96 ;
   RECT 0.0 471.96 272.84 473.67 ;
   RECT 0.0 473.67 272.84 475.38 ;
  LAYER metal4 ;
   RECT 0.0 0.0 272.84 1.71 ;
   RECT 0.0 1.71 272.84 3.42 ;
   RECT 0.0 3.42 272.84 5.13 ;
   RECT 0.0 5.13 272.84 6.84 ;
   RECT 0.0 6.84 272.84 8.55 ;
   RECT 0.0 8.55 272.84 10.26 ;
   RECT 0.0 10.26 272.84 11.97 ;
   RECT 0.0 11.97 272.84 13.68 ;
   RECT 0.0 13.68 272.84 15.39 ;
   RECT 0.0 15.39 272.84 17.1 ;
   RECT 0.0 17.1 272.84 18.81 ;
   RECT 0.0 18.81 272.84 20.52 ;
   RECT 0.0 20.52 272.84 22.23 ;
   RECT 0.0 22.23 272.84 23.94 ;
   RECT 0.0 23.94 272.84 25.65 ;
   RECT 0.0 25.65 272.84 27.36 ;
   RECT 0.0 27.36 272.84 29.07 ;
   RECT 0.0 29.07 272.84 30.78 ;
   RECT 0.0 30.78 272.84 32.49 ;
   RECT 0.0 32.49 272.84 34.2 ;
   RECT 0.0 34.2 272.84 35.91 ;
   RECT 0.0 35.91 272.84 37.62 ;
   RECT 0.0 37.62 272.84 39.33 ;
   RECT 0.0 39.33 272.84 41.04 ;
   RECT 0.0 41.04 272.84 42.75 ;
   RECT 0.0 42.75 272.84 44.46 ;
   RECT 0.0 44.46 272.84 46.17 ;
   RECT 0.0 46.17 272.84 47.88 ;
   RECT 0.0 47.88 272.84 49.59 ;
   RECT 0.0 49.59 272.84 51.3 ;
   RECT 0.0 51.3 272.84 53.01 ;
   RECT 0.0 53.01 272.84 54.72 ;
   RECT 0.0 54.72 272.84 56.43 ;
   RECT 0.0 56.43 272.84 58.14 ;
   RECT 0.0 58.14 272.84 59.85 ;
   RECT 0.0 59.85 272.84 61.56 ;
   RECT 0.0 61.56 272.84 63.27 ;
   RECT 0.0 63.27 272.84 64.98 ;
   RECT 0.0 64.98 272.84 66.69 ;
   RECT 0.0 66.69 272.84 68.4 ;
   RECT 0.0 68.4 272.84 70.11 ;
   RECT 0.0 70.11 272.84 71.82 ;
   RECT 0.0 71.82 272.84 73.53 ;
   RECT 0.0 73.53 272.84 75.24 ;
   RECT 0.0 75.24 272.84 76.95 ;
   RECT 0.0 76.95 272.84 78.66 ;
   RECT 0.0 78.66 272.84 80.37 ;
   RECT 0.0 80.37 272.84 82.08 ;
   RECT 0.0 82.08 272.84 83.79 ;
   RECT 0.0 83.79 272.84 85.5 ;
   RECT 0.0 85.5 272.84 87.21 ;
   RECT 0.0 87.21 272.84 88.92 ;
   RECT 0.0 88.92 272.84 90.63 ;
   RECT 0.0 90.63 272.84 92.34 ;
   RECT 0.0 92.34 272.84 94.05 ;
   RECT 0.0 94.05 272.84 95.76 ;
   RECT 0.0 95.76 272.84 97.47 ;
   RECT 0.0 97.47 272.84 99.18 ;
   RECT 0.0 99.18 272.84 100.89 ;
   RECT 0.0 100.89 272.84 102.6 ;
   RECT 0.0 102.6 272.84 104.31 ;
   RECT 0.0 104.31 272.84 106.02 ;
   RECT 0.0 106.02 272.84 107.73 ;
   RECT 0.0 107.73 272.84 109.44 ;
   RECT 0.0 109.44 272.84 111.15 ;
   RECT 0.0 111.15 272.84 112.86 ;
   RECT 0.0 112.86 272.84 114.57 ;
   RECT 0.0 114.57 272.84 116.28 ;
   RECT 0.0 116.28 272.84 117.99 ;
   RECT 0.0 117.99 272.84 119.7 ;
   RECT 0.0 119.7 272.84 121.41 ;
   RECT 0.0 121.41 272.84 123.12 ;
   RECT 0.0 123.12 272.84 124.83 ;
   RECT 0.0 124.83 272.84 126.54 ;
   RECT 0.0 126.54 272.84 128.25 ;
   RECT 0.0 128.25 272.84 129.96 ;
   RECT 0.0 129.96 272.84 131.67 ;
   RECT 0.0 131.67 272.84 133.38 ;
   RECT 0.0 133.38 272.84 135.09 ;
   RECT 0.0 135.09 272.84 136.8 ;
   RECT 0.0 136.8 272.84 138.51 ;
   RECT 0.0 138.51 272.84 140.22 ;
   RECT 0.0 140.22 272.84 141.93 ;
   RECT 0.0 141.93 272.84 143.64 ;
   RECT 0.0 143.64 272.84 145.35 ;
   RECT 0.0 145.35 272.84 147.06 ;
   RECT 0.0 147.06 272.84 148.77 ;
   RECT 0.0 148.77 272.84 150.48 ;
   RECT 0.0 150.48 272.84 152.19 ;
   RECT 0.0 152.19 272.84 153.9 ;
   RECT 0.0 153.9 272.84 155.61 ;
   RECT 0.0 155.61 272.84 157.32 ;
   RECT 0.0 157.32 272.84 159.03 ;
   RECT 0.0 159.03 272.84 160.74 ;
   RECT 0.0 160.74 272.84 162.45 ;
   RECT 0.0 162.45 272.84 164.16 ;
   RECT 0.0 164.16 272.84 165.87 ;
   RECT 0.0 165.87 272.84 167.58 ;
   RECT 0.0 167.58 272.84 169.29 ;
   RECT 0.0 169.29 272.84 171.0 ;
   RECT 0.0 171.0 272.84 172.71 ;
   RECT 0.0 172.71 272.84 174.42 ;
   RECT 0.0 174.42 272.84 176.13 ;
   RECT 0.0 176.13 272.84 177.84 ;
   RECT 0.0 177.84 272.84 179.55 ;
   RECT 0.0 179.55 272.84 181.26 ;
   RECT 0.0 181.26 272.84 182.97 ;
   RECT 0.0 182.97 272.84 184.68 ;
   RECT 0.0 184.68 272.84 186.39 ;
   RECT 0.0 186.39 272.84 188.1 ;
   RECT 0.0 188.1 272.84 189.81 ;
   RECT 0.0 189.81 272.84 191.52 ;
   RECT 0.0 191.52 272.84 193.23 ;
   RECT 0.0 193.23 272.84 194.94 ;
   RECT 0.0 194.94 272.84 196.65 ;
   RECT 0.0 196.65 272.84 198.36 ;
   RECT 0.0 198.36 272.84 200.07 ;
   RECT 0.0 200.07 272.84 201.78 ;
   RECT 0.0 201.78 272.84 203.49 ;
   RECT 0.0 203.49 272.84 205.2 ;
   RECT 0.0 205.2 272.84 206.91 ;
   RECT 0.0 206.91 272.84 208.62 ;
   RECT 0.0 208.62 272.84 210.33 ;
   RECT 0.0 210.33 272.84 212.04 ;
   RECT 0.0 212.04 272.84 213.75 ;
   RECT 0.0 213.75 296.02 215.46 ;
   RECT 0.0 215.46 296.02 217.17 ;
   RECT 0.0 217.17 296.02 218.88 ;
   RECT 0.0 218.88 296.02 220.59 ;
   RECT 0.0 220.59 296.02 222.3 ;
   RECT 0.0 222.3 296.02 224.01 ;
   RECT 0.0 224.01 296.02 225.72 ;
   RECT 0.0 225.72 296.02 227.43 ;
   RECT 0.0 227.43 296.02 229.14 ;
   RECT 0.0 229.14 296.02 230.85 ;
   RECT 0.0 230.85 296.02 232.56 ;
   RECT 0.0 232.56 296.02 234.27 ;
   RECT 0.0 234.27 296.02 235.98 ;
   RECT 0.0 235.98 296.02 237.69 ;
   RECT 0.0 237.69 296.02 239.4 ;
   RECT 0.0 239.4 296.02 241.11 ;
   RECT 0.0 241.11 296.02 242.82 ;
   RECT 0.0 242.82 272.84 244.53 ;
   RECT 0.0 244.53 272.84 246.24 ;
   RECT 0.0 246.24 272.84 247.95 ;
   RECT 0.0 247.95 272.84 249.66 ;
   RECT 0.0 249.66 272.84 251.37 ;
   RECT 0.0 251.37 272.84 253.08 ;
   RECT 0.0 253.08 272.84 254.79 ;
   RECT 0.0 254.79 272.84 256.5 ;
   RECT 0.0 256.5 272.84 258.21 ;
   RECT 0.0 258.21 272.84 259.92 ;
   RECT 0.0 259.92 272.84 261.63 ;
   RECT 0.0 261.63 272.84 263.34 ;
   RECT 0.0 263.34 272.84 265.05 ;
   RECT 0.0 265.05 272.84 266.76 ;
   RECT 0.0 266.76 272.84 268.47 ;
   RECT 0.0 268.47 272.84 270.18 ;
   RECT 0.0 270.18 272.84 271.89 ;
   RECT 0.0 271.89 272.84 273.6 ;
   RECT 0.0 273.6 272.84 275.31 ;
   RECT 0.0 275.31 272.84 277.02 ;
   RECT 0.0 277.02 272.84 278.73 ;
   RECT 0.0 278.73 272.84 280.44 ;
   RECT 0.0 280.44 272.84 282.15 ;
   RECT 0.0 282.15 272.84 283.86 ;
   RECT 0.0 283.86 272.84 285.57 ;
   RECT 0.0 285.57 272.84 287.28 ;
   RECT 0.0 287.28 272.84 288.99 ;
   RECT 0.0 288.99 272.84 290.7 ;
   RECT 0.0 290.7 272.84 292.41 ;
   RECT 0.0 292.41 272.84 294.12 ;
   RECT 0.0 294.12 272.84 295.83 ;
   RECT 0.0 295.83 272.84 297.54 ;
   RECT 0.0 297.54 272.84 299.25 ;
   RECT 0.0 299.25 272.84 300.96 ;
   RECT 0.0 300.96 272.84 302.67 ;
   RECT 0.0 302.67 272.84 304.38 ;
   RECT 0.0 304.38 272.84 306.09 ;
   RECT 0.0 306.09 272.84 307.8 ;
   RECT 0.0 307.8 272.84 309.51 ;
   RECT 0.0 309.51 272.84 311.22 ;
   RECT 0.0 311.22 272.84 312.93 ;
   RECT 0.0 312.93 272.84 314.64 ;
   RECT 0.0 314.64 272.84 316.35 ;
   RECT 0.0 316.35 272.84 318.06 ;
   RECT 0.0 318.06 272.84 319.77 ;
   RECT 0.0 319.77 272.84 321.48 ;
   RECT 0.0 321.48 272.84 323.19 ;
   RECT 0.0 323.19 272.84 324.9 ;
   RECT 0.0 324.9 272.84 326.61 ;
   RECT 0.0 326.61 272.84 328.32 ;
   RECT 0.0 328.32 272.84 330.03 ;
   RECT 0.0 330.03 272.84 331.74 ;
   RECT 0.0 331.74 272.84 333.45 ;
   RECT 0.0 333.45 272.84 335.16 ;
   RECT 0.0 335.16 272.84 336.87 ;
   RECT 0.0 336.87 272.84 338.58 ;
   RECT 0.0 338.58 272.84 340.29 ;
   RECT 0.0 340.29 272.84 342.0 ;
   RECT 0.0 342.0 272.84 343.71 ;
   RECT 0.0 343.71 272.84 345.42 ;
   RECT 0.0 345.42 272.84 347.13 ;
   RECT 0.0 347.13 272.84 348.84 ;
   RECT 0.0 348.84 272.84 350.55 ;
   RECT 0.0 350.55 272.84 352.26 ;
   RECT 0.0 352.26 272.84 353.97 ;
   RECT 0.0 353.97 272.84 355.68 ;
   RECT 0.0 355.68 272.84 357.39 ;
   RECT 0.0 357.39 272.84 359.1 ;
   RECT 0.0 359.1 272.84 360.81 ;
   RECT 0.0 360.81 272.84 362.52 ;
   RECT 0.0 362.52 272.84 364.23 ;
   RECT 0.0 364.23 272.84 365.94 ;
   RECT 0.0 365.94 272.84 367.65 ;
   RECT 0.0 367.65 272.84 369.36 ;
   RECT 0.0 369.36 272.84 371.07 ;
   RECT 0.0 371.07 272.84 372.78 ;
   RECT 0.0 372.78 272.84 374.49 ;
   RECT 0.0 374.49 272.84 376.2 ;
   RECT 0.0 376.2 272.84 377.91 ;
   RECT 0.0 377.91 272.84 379.62 ;
   RECT 0.0 379.62 272.84 381.33 ;
   RECT 0.0 381.33 272.84 383.04 ;
   RECT 0.0 383.04 272.84 384.75 ;
   RECT 0.0 384.75 272.84 386.46 ;
   RECT 0.0 386.46 272.84 388.17 ;
   RECT 0.0 388.17 272.84 389.88 ;
   RECT 0.0 389.88 272.84 391.59 ;
   RECT 0.0 391.59 272.84 393.3 ;
   RECT 0.0 393.3 272.84 395.01 ;
   RECT 0.0 395.01 272.84 396.72 ;
   RECT 0.0 396.72 272.84 398.43 ;
   RECT 0.0 398.43 272.84 400.14 ;
   RECT 0.0 400.14 272.84 401.85 ;
   RECT 0.0 401.85 272.84 403.56 ;
   RECT 0.0 403.56 272.84 405.27 ;
   RECT 0.0 405.27 272.84 406.98 ;
   RECT 0.0 406.98 272.84 408.69 ;
   RECT 0.0 408.69 272.84 410.4 ;
   RECT 0.0 410.4 272.84 412.11 ;
   RECT 0.0 412.11 272.84 413.82 ;
   RECT 0.0 413.82 272.84 415.53 ;
   RECT 0.0 415.53 272.84 417.24 ;
   RECT 0.0 417.24 272.84 418.95 ;
   RECT 0.0 418.95 272.84 420.66 ;
   RECT 0.0 420.66 272.84 422.37 ;
   RECT 0.0 422.37 272.84 424.08 ;
   RECT 0.0 424.08 272.84 425.79 ;
   RECT 0.0 425.79 272.84 427.5 ;
   RECT 0.0 427.5 272.84 429.21 ;
   RECT 0.0 429.21 272.84 430.92 ;
   RECT 0.0 430.92 272.84 432.63 ;
   RECT 0.0 432.63 272.84 434.34 ;
   RECT 0.0 434.34 272.84 436.05 ;
   RECT 0.0 436.05 272.84 437.76 ;
   RECT 0.0 437.76 272.84 439.47 ;
   RECT 0.0 439.47 272.84 441.18 ;
   RECT 0.0 441.18 272.84 442.89 ;
   RECT 0.0 442.89 272.84 444.6 ;
   RECT 0.0 444.6 272.84 446.31 ;
   RECT 0.0 446.31 272.84 448.02 ;
   RECT 0.0 448.02 272.84 449.73 ;
   RECT 0.0 449.73 272.84 451.44 ;
   RECT 0.0 451.44 272.84 453.15 ;
   RECT 0.0 453.15 272.84 454.86 ;
   RECT 0.0 454.86 272.84 456.57 ;
   RECT 0.0 456.57 272.84 458.28 ;
   RECT 0.0 458.28 272.84 459.99 ;
   RECT 0.0 459.99 272.84 461.7 ;
   RECT 0.0 461.7 272.84 463.41 ;
   RECT 0.0 463.41 272.84 465.12 ;
   RECT 0.0 465.12 272.84 466.83 ;
   RECT 0.0 466.83 272.84 468.54 ;
   RECT 0.0 468.54 272.84 470.25 ;
   RECT 0.0 470.25 272.84 471.96 ;
   RECT 0.0 471.96 272.84 473.67 ;
   RECT 0.0 473.67 272.84 475.38 ;
 END
END block_779x2502_158

MACRO block_341x369_80
 CLASS BLOCK ;
 FOREIGN block_341x369_80 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 129.58 BY 70.11 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 20.235 126.445 20.805 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 26.695 126.445 27.265 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 6.935 3.325 7.505 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 9.215 3.325 9.785 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 10.735 3.325 11.305 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 13.015 3.325 13.585 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 13.395 4.085 13.965 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 13.775 3.325 14.345 ;
  END
 END o7
 PIN o8
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 15.295 3.325 15.865 ;
  END
 END o8
 PIN o9
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 16.055 3.325 16.625 ;
  END
 END o9
 PIN o10
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 16.815 3.325 17.385 ;
  END
 END o10
 PIN o11
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 12.635 4.085 13.205 ;
  END
 END o11
 PIN o12
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 19.855 3.325 20.425 ;
  END
 END o12
 PIN o13
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 20.615 3.325 21.185 ;
  END
 END o13
 PIN o14
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 21.375 3.325 21.945 ;
  END
 END o14
 PIN o15
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 22.135 3.325 22.705 ;
  END
 END o15
 PIN o16
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 22.895 3.325 23.465 ;
  END
 END o16
 PIN o17
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 18.335 3.325 18.905 ;
  END
 END o17
 PIN o18
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 25.935 3.325 26.505 ;
  END
 END o18
 PIN o19
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 26.695 3.325 27.265 ;
  END
 END o19
 PIN o20
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 27.455 3.325 28.025 ;
  END
 END o20
 PIN o21
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 28.975 3.325 29.545 ;
  END
 END o21
 PIN o22
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 29.735 3.325 30.305 ;
  END
 END o22
 PIN o23
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 25.175 3.325 25.745 ;
  END
 END o23
 PIN o24
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 32.015 3.325 32.585 ;
  END
 END o24
 PIN o25
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 33.535 3.325 34.105 ;
  END
 END o25
 PIN o26
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 34.295 3.325 34.865 ;
  END
 END o26
 PIN o27
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 35.055 3.325 35.625 ;
  END
 END o27
 PIN o28
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 35.815 3.325 36.385 ;
  END
 END o28
 PIN o29
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 31.255 3.325 31.825 ;
  END
 END o29
 PIN o30
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 38.095 126.445 38.665 ;
  END
 END o30
 PIN o31
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 38.855 126.445 39.425 ;
  END
 END o31
 PIN o32
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 39.615 126.445 40.185 ;
  END
 END o32
 PIN o33
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 42.655 126.445 43.225 ;
  END
 END o33
 PIN o34
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 29.735 126.445 30.305 ;
  END
 END o34
 PIN o35
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 21.755 126.445 22.325 ;
  END
 END o35
 PIN o36
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 31.255 126.445 31.825 ;
  END
 END o36
 PIN o37
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 32.015 126.445 32.585 ;
  END
 END o37
 PIN o38
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 33.535 126.445 34.105 ;
  END
 END o38
 PIN o39
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 34.295 126.445 34.865 ;
  END
 END o39
 PIN o40
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 35.055 126.445 35.625 ;
  END
 END o40
 PIN o41
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 30.495 126.445 31.065 ;
  END
 END o41
 PIN o42
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 28.975 126.445 29.545 ;
  END
 END o42
 PIN o43
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 41.135 3.325 41.705 ;
  END
 END o43
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 35.815 126.445 36.385 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 43.035 125.685 43.605 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 32.395 125.685 32.965 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 35.435 125.685 36.005 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 36.955 126.445 37.525 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 36.575 125.685 37.145 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 33.915 125.685 34.485 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 30.115 125.685 30.685 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 40.375 3.325 40.945 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 8.455 3.325 9.025 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 25.935 126.445 26.505 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 25.175 126.445 25.745 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 24.415 126.445 24.985 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 34.675 125.685 35.245 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 30.875 125.685 31.445 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 40.755 126.445 41.325 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 27.455 126.445 28.025 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 38.475 125.685 39.045 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 39.995 125.685 40.565 ;
  END
 END i18
 PIN i19
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 39.235 125.685 39.805 ;
  END
 END i19
 PIN i20
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 124.355 40.375 124.925 40.945 ;
  END
 END i20
 PIN i21
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 8.455 126.445 9.025 ;
  END
 END i21
 PIN i22
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 9.215 126.445 9.785 ;
  END
 END i22
 PIN i23
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 10.735 126.445 11.305 ;
  END
 END i23
 PIN i24
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 11.495 126.445 12.065 ;
  END
 END i24
 PIN i25
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 12.255 126.445 12.825 ;
  END
 END i25
 PIN i26
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 13.015 126.445 13.585 ;
  END
 END i26
 PIN i27
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 8.075 125.685 8.645 ;
  END
 END i27
 PIN i28
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 7.695 126.445 8.265 ;
  END
 END i28
 PIN i29
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 7.315 125.685 7.885 ;
  END
 END i29
 PIN i30
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 6.935 126.445 7.505 ;
  END
 END i30
 PIN i31
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 6.555 125.685 7.125 ;
  END
 END i31
 PIN i32
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 13.775 126.445 14.345 ;
  END
 END i32
 PIN i33
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 15.295 126.445 15.865 ;
  END
 END i33
 PIN i34
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 16.055 126.445 16.625 ;
  END
 END i34
 PIN i35
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 16.815 126.445 17.385 ;
  END
 END i35
 OBS
  LAYER metal1 ;
   RECT 0 0 129.58 70.11 ;
  LAYER via1 ;
   RECT 0 0 129.58 70.11 ;
  LAYER metal2 ;
   RECT 0 0 129.58 70.11 ;
  LAYER via2 ;
   RECT 0 0 129.58 70.11 ;
  LAYER metal3 ;
   RECT 0 0 129.58 70.11 ;
  LAYER via3 ;
   RECT 0 0 129.58 70.11 ;
  LAYER metal4 ;
   RECT 0 0 129.58 70.11 ;
 END
END block_341x369_80

MACRO block_1024x2502_161
 CLASS BLOCK ;
 FOREIGN block_1024x2502_161 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 389.12 BY 475.38 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 8.455 362.805 9.025 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 24.795 362.805 25.365 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 190.095 362.805 190.665 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 206.435 362.805 207.005 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 222.775 362.805 223.345 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 267.235 362.805 267.805 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 283.575 362.805 284.145 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 299.915 362.805 300.485 ;
  END
 END o7
 PIN o8
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 316.255 362.805 316.825 ;
  END
 END o8
 PIN o9
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 332.595 362.805 333.165 ;
  END
 END o9
 PIN o10
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 348.935 362.805 349.505 ;
  END
 END o10
 PIN o11
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 383.515 362.805 384.085 ;
  END
 END o11
 PIN o12
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 41.135 362.805 41.705 ;
  END
 END o12
 PIN o13
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 399.855 362.805 400.425 ;
  END
 END o13
 PIN o14
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 416.195 362.805 416.765 ;
  END
 END o14
 PIN o15
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 432.535 362.805 433.105 ;
  END
 END o15
 PIN o16
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 448.875 362.805 449.445 ;
  END
 END o16
 PIN o17
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 465.215 362.805 465.785 ;
  END
 END o17
 PIN o18
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 57.475 362.805 58.045 ;
  END
 END o18
 PIN o19
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 73.815 362.805 74.385 ;
  END
 END o19
 PIN o20
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 90.155 362.805 90.725 ;
  END
 END o20
 PIN o21
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 106.495 362.805 107.065 ;
  END
 END o21
 PIN o22
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 141.075 362.805 141.645 ;
  END
 END o22
 PIN o23
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 157.415 362.805 157.985 ;
  END
 END o23
 PIN o24
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 173.755 362.805 174.325 ;
  END
 END o24
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 385.415 233.795 385.985 234.365 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 385.415 250.895 385.985 251.465 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 385.415 239.115 385.985 239.685 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 385.415 243.485 385.985 244.055 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 385.415 246.335 385.985 246.905 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 384.655 234.175 385.225 234.745 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 384.655 233.415 385.225 233.985 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 385.415 233.035 385.985 233.605 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 385.415 242.725 385.985 243.295 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 385.415 255.835 385.985 256.405 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 384.655 250.515 385.225 251.085 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 385.415 247.285 385.985 247.855 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 385.415 254.695 385.985 255.265 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 385.415 250.135 385.985 250.705 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 385.415 252.225 385.985 252.795 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 384.655 255.075 385.225 255.645 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 384.655 256.215 385.225 256.785 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 374.395 232.655 374.965 233.225 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 374.395 245.955 374.965 246.525 ;
  END
 END i18
 PIN i19
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 6.745 362.805 7.315 ;
  END
 END i19
 PIN i20
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 23.085 362.805 23.655 ;
  END
 END i20
 PIN i21
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 188.385 362.805 188.955 ;
  END
 END i21
 PIN i22
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 204.725 362.805 205.295 ;
  END
 END i22
 PIN i23
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 221.065 362.805 221.635 ;
  END
 END i23
 PIN i24
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 268.945 362.805 269.515 ;
  END
 END i24
 PIN i25
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 285.285 362.805 285.855 ;
  END
 END i25
 PIN i26
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 301.625 362.805 302.195 ;
  END
 END i26
 PIN i27
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 317.965 362.805 318.535 ;
  END
 END i27
 PIN i28
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 334.305 362.805 334.875 ;
  END
 END i28
 PIN i29
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 350.645 362.805 351.215 ;
  END
 END i29
 PIN i30
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 385.225 362.805 385.795 ;
  END
 END i30
 PIN i31
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 39.425 362.805 39.995 ;
  END
 END i31
 PIN i32
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 401.565 362.805 402.135 ;
  END
 END i32
 PIN i33
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 417.905 362.805 418.475 ;
  END
 END i33
 PIN i34
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 434.245 362.805 434.815 ;
  END
 END i34
 PIN i35
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 450.585 362.805 451.155 ;
  END
 END i35
 PIN i36
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 466.925 362.805 467.495 ;
  END
 END i36
 PIN i37
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 55.765 362.805 56.335 ;
  END
 END i37
 PIN i38
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 72.105 362.805 72.675 ;
  END
 END i38
 PIN i39
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 88.445 362.805 89.015 ;
  END
 END i39
 PIN i40
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 104.785 362.805 105.355 ;
  END
 END i40
 PIN i41
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 139.365 362.805 139.935 ;
  END
 END i41
 PIN i42
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 155.705 362.805 156.275 ;
  END
 END i42
 PIN i43
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 172.045 362.805 172.615 ;
  END
 END i43
 PIN i44
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 361.475 90.725 362.045 91.295 ;
  END
 END i44
 PIN i45
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 94.715 362.805 95.285 ;
  END
 END i45
 PIN i46
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 98.895 362.805 99.465 ;
  END
 END i46
 PIN i47
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 78.375 362.805 78.945 ;
  END
 END i47
 PIN i48
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 82.555 362.805 83.125 ;
  END
 END i48
 PIN i49
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 361.475 157.985 362.045 158.555 ;
  END
 END i49
 PIN i50
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 161.975 362.805 162.545 ;
  END
 END i50
 PIN i51
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 166.155 362.805 166.725 ;
  END
 END i51
 PIN i52
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 170.145 362.805 170.715 ;
  END
 END i52
 PIN i53
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 361.475 174.325 362.045 174.895 ;
  END
 END i53
 PIN i54
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 361.475 332.025 362.045 332.595 ;
  END
 END i54
 PIN i55
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 328.035 362.805 328.605 ;
  END
 END i55
 PIN i56
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 323.855 362.805 324.425 ;
  END
 END i56
 PIN i57
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 319.865 362.805 320.435 ;
  END
 END i57
 PIN i58
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 361.475 315.685 362.045 316.255 ;
  END
 END i58
 PIN i59
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 361.475 399.285 362.045 399.855 ;
  END
 END i59
 PIN i60
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 395.295 362.805 395.865 ;
  END
 END i60
 PIN i61
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 391.115 362.805 391.685 ;
  END
 END i61
 PIN i62
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 411.635 362.805 412.205 ;
  END
 END i62
 PIN i63
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 407.455 362.805 408.025 ;
  END
 END i63
 PIN i64
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 86.545 362.805 87.115 ;
  END
 END i64
 PIN i65
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 153.805 362.805 154.375 ;
  END
 END i65
 PIN i66
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 336.205 362.805 336.775 ;
  END
 END i66
 PIN i67
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 362.235 403.465 362.805 404.035 ;
  END
 END i67
 PIN i68
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 370.595 232.655 371.165 233.225 ;
  END
 END i68
 PIN i69
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 370.595 245.955 371.165 246.525 ;
  END
 END i69
 PIN i70
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 361.475 7.315 362.045 7.885 ;
  END
 END i70
 PIN i71
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 361.475 23.655 362.045 24.225 ;
  END
 END i71
 PIN i72
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 361.475 188.955 362.045 189.525 ;
  END
 END i72
 PIN i73
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 361.475 205.295 362.045 205.865 ;
  END
 END i73
 PIN i74
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 361.475 221.635 362.045 222.205 ;
  END
 END i74
 PIN i75
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 361.475 268.375 362.045 268.945 ;
  END
 END i75
 PIN i76
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 361.475 284.715 362.045 285.285 ;
  END
 END i76
 PIN i77
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 361.475 301.055 362.045 301.625 ;
  END
 END i77
 PIN i78
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 361.475 317.395 362.045 317.965 ;
  END
 END i78
 PIN i79
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 361.475 333.735 362.045 334.305 ;
  END
 END i79
 PIN i80
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 361.475 350.075 362.045 350.645 ;
  END
 END i80
 PIN i81
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 361.475 384.655 362.045 385.225 ;
  END
 END i81
 PIN i82
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 361.475 39.995 362.045 40.565 ;
  END
 END i82
 PIN i83
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 361.475 400.995 362.045 401.565 ;
  END
 END i83
 PIN i84
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 361.475 417.335 362.045 417.905 ;
  END
 END i84
 PIN i85
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 361.475 433.675 362.045 434.245 ;
  END
 END i85
 PIN i86
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 361.475 450.015 362.045 450.585 ;
  END
 END i86
 PIN i87
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 361.475 466.355 362.045 466.925 ;
  END
 END i87
 PIN i88
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 361.475 56.335 362.045 56.905 ;
  END
 END i88
 PIN i89
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 361.475 72.675 362.045 73.245 ;
  END
 END i89
 PIN i90
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 361.475 89.015 362.045 89.585 ;
  END
 END i90
 PIN i91
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 361.475 105.355 362.045 105.925 ;
  END
 END i91
 PIN i92
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 361.475 139.935 362.045 140.505 ;
  END
 END i92
 PIN i93
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 361.475 156.275 362.045 156.845 ;
  END
 END i93
 PIN i94
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 361.475 172.615 362.045 173.185 ;
  END
 END i94
 PIN i95
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 385.415 240.255 385.985 240.825 ;
  END
 END i95
 PIN i96
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 384.655 240.635 385.225 241.205 ;
  END
 END i96
 PIN i97
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 360.715 7.885 361.285 8.455 ;
  END
 END i97
 PIN i98
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 360.715 24.225 361.285 24.795 ;
  END
 END i98
 PIN i99
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 360.715 189.525 361.285 190.095 ;
  END
 END i99
 PIN i100
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 360.715 205.865 361.285 206.435 ;
  END
 END i100
 PIN i101
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 360.715 222.205 361.285 222.775 ;
  END
 END i101
 PIN i102
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 360.715 267.805 361.285 268.375 ;
  END
 END i102
 PIN i103
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 360.715 284.145 361.285 284.715 ;
  END
 END i103
 PIN i104
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 360.715 300.485 361.285 301.055 ;
  END
 END i104
 PIN i105
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 360.715 316.825 361.285 317.395 ;
  END
 END i105
 PIN i106
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 360.715 333.165 361.285 333.735 ;
  END
 END i106
 PIN i107
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 360.715 349.505 361.285 350.075 ;
  END
 END i107
 PIN i108
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 360.715 384.085 361.285 384.655 ;
  END
 END i108
 PIN i109
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 360.715 40.565 361.285 41.135 ;
  END
 END i109
 PIN i110
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 360.715 400.425 361.285 400.995 ;
  END
 END i110
 PIN i111
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 360.715 416.765 361.285 417.335 ;
  END
 END i111
 PIN i112
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 360.715 433.105 361.285 433.675 ;
  END
 END i112
 PIN i113
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 360.715 449.445 361.285 450.015 ;
  END
 END i113
 PIN i114
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 360.715 465.785 361.285 466.355 ;
  END
 END i114
 PIN i115
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 360.715 56.905 361.285 57.475 ;
  END
 END i115
 PIN i116
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 360.715 73.245 361.285 73.815 ;
  END
 END i116
 PIN i117
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 360.715 89.585 361.285 90.155 ;
  END
 END i117
 PIN i118
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 360.715 105.925 361.285 106.495 ;
  END
 END i118
 PIN i119
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 360.715 140.505 361.285 141.075 ;
  END
 END i119
 PIN i120
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 360.715 156.845 361.285 157.415 ;
  END
 END i120
 PIN i121
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 360.715 173.185 361.285 173.755 ;
  END
 END i121
 PIN i122
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 384.275 232.655 384.845 233.225 ;
  END
 END i122
 PIN i123
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 383.135 232.655 383.705 233.225 ;
  END
 END i123
 PIN i124
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 381.615 232.655 382.185 233.225 ;
  END
 END i124
 PIN i125
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 379.715 232.655 380.285 233.225 ;
  END
 END i125
 PIN i126
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 378.575 232.655 379.145 233.225 ;
  END
 END i126
 PIN i127
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 376.675 232.655 377.245 233.225 ;
  END
 END i127
 PIN i128
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 375.535 232.655 376.105 233.225 ;
  END
 END i128
 PIN i129
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 384.275 245.955 384.845 246.525 ;
  END
 END i129
 PIN i130
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 383.135 245.955 383.705 246.525 ;
  END
 END i130
 PIN i131
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 381.615 245.955 382.185 246.525 ;
  END
 END i131
 PIN i132
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 379.715 245.955 380.285 246.525 ;
  END
 END i132
 PIN i133
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 378.575 245.955 379.145 246.525 ;
  END
 END i133
 PIN i134
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 376.675 245.955 377.245 246.525 ;
  END
 END i134
 PIN i135
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 375.535 245.955 376.105 246.525 ;
  END
 END i135
 OBS
  LAYER metal1 ;
   RECT 0.0 0.0 365.94 1.71 ;
   RECT 0.0 1.71 365.94 3.42 ;
   RECT 0.0 3.42 365.94 5.13 ;
   RECT 0.0 5.13 365.94 6.84 ;
   RECT 0.0 6.84 365.94 8.55 ;
   RECT 0.0 8.55 365.94 10.26 ;
   RECT 0.0 10.26 365.94 11.97 ;
   RECT 0.0 11.97 365.94 13.68 ;
   RECT 0.0 13.68 365.94 15.39 ;
   RECT 0.0 15.39 365.94 17.1 ;
   RECT 0.0 17.1 365.94 18.81 ;
   RECT 0.0 18.81 365.94 20.52 ;
   RECT 0.0 20.52 365.94 22.23 ;
   RECT 0.0 22.23 365.94 23.94 ;
   RECT 0.0 23.94 365.94 25.65 ;
   RECT 0.0 25.65 365.94 27.36 ;
   RECT 0.0 27.36 365.94 29.07 ;
   RECT 0.0 29.07 365.94 30.78 ;
   RECT 0.0 30.78 365.94 32.49 ;
   RECT 0.0 32.49 365.94 34.2 ;
   RECT 0.0 34.2 365.94 35.91 ;
   RECT 0.0 35.91 365.94 37.62 ;
   RECT 0.0 37.62 365.94 39.33 ;
   RECT 0.0 39.33 365.94 41.04 ;
   RECT 0.0 41.04 365.94 42.75 ;
   RECT 0.0 42.75 365.94 44.46 ;
   RECT 0.0 44.46 365.94 46.17 ;
   RECT 0.0 46.17 365.94 47.88 ;
   RECT 0.0 47.88 365.94 49.59 ;
   RECT 0.0 49.59 365.94 51.3 ;
   RECT 0.0 51.3 365.94 53.01 ;
   RECT 0.0 53.01 365.94 54.72 ;
   RECT 0.0 54.72 365.94 56.43 ;
   RECT 0.0 56.43 365.94 58.14 ;
   RECT 0.0 58.14 365.94 59.85 ;
   RECT 0.0 59.85 365.94 61.56 ;
   RECT 0.0 61.56 365.94 63.27 ;
   RECT 0.0 63.27 365.94 64.98 ;
   RECT 0.0 64.98 365.94 66.69 ;
   RECT 0.0 66.69 365.94 68.4 ;
   RECT 0.0 68.4 365.94 70.11 ;
   RECT 0.0 70.11 365.94 71.82 ;
   RECT 0.0 71.82 365.94 73.53 ;
   RECT 0.0 73.53 365.94 75.24 ;
   RECT 0.0 75.24 365.94 76.95 ;
   RECT 0.0 76.95 365.94 78.66 ;
   RECT 0.0 78.66 365.94 80.37 ;
   RECT 0.0 80.37 365.94 82.08 ;
   RECT 0.0 82.08 365.94 83.79 ;
   RECT 0.0 83.79 365.94 85.5 ;
   RECT 0.0 85.5 365.94 87.21 ;
   RECT 0.0 87.21 365.94 88.92 ;
   RECT 0.0 88.92 365.94 90.63 ;
   RECT 0.0 90.63 365.94 92.34 ;
   RECT 0.0 92.34 365.94 94.05 ;
   RECT 0.0 94.05 365.94 95.76 ;
   RECT 0.0 95.76 365.94 97.47 ;
   RECT 0.0 97.47 365.94 99.18 ;
   RECT 0.0 99.18 365.94 100.89 ;
   RECT 0.0 100.89 365.94 102.6 ;
   RECT 0.0 102.6 365.94 104.31 ;
   RECT 0.0 104.31 365.94 106.02 ;
   RECT 0.0 106.02 365.94 107.73 ;
   RECT 0.0 107.73 365.94 109.44 ;
   RECT 0.0 109.44 365.94 111.15 ;
   RECT 0.0 111.15 365.94 112.86 ;
   RECT 0.0 112.86 365.94 114.57 ;
   RECT 0.0 114.57 365.94 116.28 ;
   RECT 0.0 116.28 365.94 117.99 ;
   RECT 0.0 117.99 365.94 119.7 ;
   RECT 0.0 119.7 365.94 121.41 ;
   RECT 0.0 121.41 365.94 123.12 ;
   RECT 0.0 123.12 365.94 124.83 ;
   RECT 0.0 124.83 365.94 126.54 ;
   RECT 0.0 126.54 365.94 128.25 ;
   RECT 0.0 128.25 365.94 129.96 ;
   RECT 0.0 129.96 365.94 131.67 ;
   RECT 0.0 131.67 365.94 133.38 ;
   RECT 0.0 133.38 365.94 135.09 ;
   RECT 0.0 135.09 365.94 136.8 ;
   RECT 0.0 136.8 365.94 138.51 ;
   RECT 0.0 138.51 365.94 140.22 ;
   RECT 0.0 140.22 365.94 141.93 ;
   RECT 0.0 141.93 365.94 143.64 ;
   RECT 0.0 143.64 365.94 145.35 ;
   RECT 0.0 145.35 365.94 147.06 ;
   RECT 0.0 147.06 365.94 148.77 ;
   RECT 0.0 148.77 365.94 150.48 ;
   RECT 0.0 150.48 365.94 152.19 ;
   RECT 0.0 152.19 365.94 153.9 ;
   RECT 0.0 153.9 365.94 155.61 ;
   RECT 0.0 155.61 365.94 157.32 ;
   RECT 0.0 157.32 365.94 159.03 ;
   RECT 0.0 159.03 365.94 160.74 ;
   RECT 0.0 160.74 365.94 162.45 ;
   RECT 0.0 162.45 365.94 164.16 ;
   RECT 0.0 164.16 365.94 165.87 ;
   RECT 0.0 165.87 365.94 167.58 ;
   RECT 0.0 167.58 365.94 169.29 ;
   RECT 0.0 169.29 365.94 171.0 ;
   RECT 0.0 171.0 365.94 172.71 ;
   RECT 0.0 172.71 365.94 174.42 ;
   RECT 0.0 174.42 365.94 176.13 ;
   RECT 0.0 176.13 365.94 177.84 ;
   RECT 0.0 177.84 365.94 179.55 ;
   RECT 0.0 179.55 365.94 181.26 ;
   RECT 0.0 181.26 365.94 182.97 ;
   RECT 0.0 182.97 365.94 184.68 ;
   RECT 0.0 184.68 365.94 186.39 ;
   RECT 0.0 186.39 365.94 188.1 ;
   RECT 0.0 188.1 365.94 189.81 ;
   RECT 0.0 189.81 365.94 191.52 ;
   RECT 0.0 191.52 365.94 193.23 ;
   RECT 0.0 193.23 365.94 194.94 ;
   RECT 0.0 194.94 365.94 196.65 ;
   RECT 0.0 196.65 365.94 198.36 ;
   RECT 0.0 198.36 365.94 200.07 ;
   RECT 0.0 200.07 365.94 201.78 ;
   RECT 0.0 201.78 365.94 203.49 ;
   RECT 0.0 203.49 365.94 205.2 ;
   RECT 0.0 205.2 365.94 206.91 ;
   RECT 0.0 206.91 365.94 208.62 ;
   RECT 0.0 208.62 365.94 210.33 ;
   RECT 0.0 210.33 365.94 212.04 ;
   RECT 0.0 212.04 365.94 213.75 ;
   RECT 0.0 213.75 365.94 215.46 ;
   RECT 0.0 215.46 365.94 217.17 ;
   RECT 0.0 217.17 365.94 218.88 ;
   RECT 0.0 218.88 365.94 220.59 ;
   RECT 0.0 220.59 365.94 222.3 ;
   RECT 0.0 222.3 365.94 224.01 ;
   RECT 0.0 224.01 365.94 225.72 ;
   RECT 0.0 225.72 365.94 227.43 ;
   RECT 0.0 227.43 365.94 229.14 ;
   RECT 0.0 229.14 365.94 230.85 ;
   RECT 0.0 230.85 389.12 232.56 ;
   RECT 0.0 232.56 389.12 234.27 ;
   RECT 0.0 234.27 389.12 235.98 ;
   RECT 0.0 235.98 389.12 237.69 ;
   RECT 0.0 237.69 389.12 239.4 ;
   RECT 0.0 239.4 389.12 241.11 ;
   RECT 0.0 241.11 389.12 242.82 ;
   RECT 0.0 242.82 389.12 244.53 ;
   RECT 0.0 244.53 389.12 246.24 ;
   RECT 0.0 246.24 389.12 247.95 ;
   RECT 0.0 247.95 389.12 249.66 ;
   RECT 0.0 249.66 389.12 251.37 ;
   RECT 0.0 251.37 389.12 253.08 ;
   RECT 0.0 253.08 389.12 254.79 ;
   RECT 0.0 254.79 389.12 256.5 ;
   RECT 0.0 256.5 389.12 258.21 ;
   RECT 0.0 258.21 389.12 259.92 ;
   RECT 0.0 259.92 365.94 261.63 ;
   RECT 0.0 261.63 365.94 263.34 ;
   RECT 0.0 263.34 365.94 265.05 ;
   RECT 0.0 265.05 365.94 266.76 ;
   RECT 0.0 266.76 365.94 268.47 ;
   RECT 0.0 268.47 365.94 270.18 ;
   RECT 0.0 270.18 365.94 271.89 ;
   RECT 0.0 271.89 365.94 273.6 ;
   RECT 0.0 273.6 365.94 275.31 ;
   RECT 0.0 275.31 365.94 277.02 ;
   RECT 0.0 277.02 365.94 278.73 ;
   RECT 0.0 278.73 365.94 280.44 ;
   RECT 0.0 280.44 365.94 282.15 ;
   RECT 0.0 282.15 365.94 283.86 ;
   RECT 0.0 283.86 365.94 285.57 ;
   RECT 0.0 285.57 365.94 287.28 ;
   RECT 0.0 287.28 365.94 288.99 ;
   RECT 0.0 288.99 365.94 290.7 ;
   RECT 0.0 290.7 365.94 292.41 ;
   RECT 0.0 292.41 365.94 294.12 ;
   RECT 0.0 294.12 365.94 295.83 ;
   RECT 0.0 295.83 365.94 297.54 ;
   RECT 0.0 297.54 365.94 299.25 ;
   RECT 0.0 299.25 365.94 300.96 ;
   RECT 0.0 300.96 365.94 302.67 ;
   RECT 0.0 302.67 365.94 304.38 ;
   RECT 0.0 304.38 365.94 306.09 ;
   RECT 0.0 306.09 365.94 307.8 ;
   RECT 0.0 307.8 365.94 309.51 ;
   RECT 0.0 309.51 365.94 311.22 ;
   RECT 0.0 311.22 365.94 312.93 ;
   RECT 0.0 312.93 365.94 314.64 ;
   RECT 0.0 314.64 365.94 316.35 ;
   RECT 0.0 316.35 365.94 318.06 ;
   RECT 0.0 318.06 365.94 319.77 ;
   RECT 0.0 319.77 365.94 321.48 ;
   RECT 0.0 321.48 365.94 323.19 ;
   RECT 0.0 323.19 365.94 324.9 ;
   RECT 0.0 324.9 365.94 326.61 ;
   RECT 0.0 326.61 365.94 328.32 ;
   RECT 0.0 328.32 365.94 330.03 ;
   RECT 0.0 330.03 365.94 331.74 ;
   RECT 0.0 331.74 365.94 333.45 ;
   RECT 0.0 333.45 365.94 335.16 ;
   RECT 0.0 335.16 365.94 336.87 ;
   RECT 0.0 336.87 365.94 338.58 ;
   RECT 0.0 338.58 365.94 340.29 ;
   RECT 0.0 340.29 365.94 342.0 ;
   RECT 0.0 342.0 365.94 343.71 ;
   RECT 0.0 343.71 365.94 345.42 ;
   RECT 0.0 345.42 365.94 347.13 ;
   RECT 0.0 347.13 365.94 348.84 ;
   RECT 0.0 348.84 365.94 350.55 ;
   RECT 0.0 350.55 365.94 352.26 ;
   RECT 0.0 352.26 365.94 353.97 ;
   RECT 0.0 353.97 365.94 355.68 ;
   RECT 0.0 355.68 365.94 357.39 ;
   RECT 0.0 357.39 365.94 359.1 ;
   RECT 0.0 359.1 365.94 360.81 ;
   RECT 0.0 360.81 365.94 362.52 ;
   RECT 0.0 362.52 365.94 364.23 ;
   RECT 0.0 364.23 365.94 365.94 ;
   RECT 0.0 365.94 365.94 367.65 ;
   RECT 0.0 367.65 365.94 369.36 ;
   RECT 0.0 369.36 365.94 371.07 ;
   RECT 0.0 371.07 365.94 372.78 ;
   RECT 0.0 372.78 365.94 374.49 ;
   RECT 0.0 374.49 365.94 376.2 ;
   RECT 0.0 376.2 365.94 377.91 ;
   RECT 0.0 377.91 365.94 379.62 ;
   RECT 0.0 379.62 365.94 381.33 ;
   RECT 0.0 381.33 365.94 383.04 ;
   RECT 0.0 383.04 365.94 384.75 ;
   RECT 0.0 384.75 365.94 386.46 ;
   RECT 0.0 386.46 365.94 388.17 ;
   RECT 0.0 388.17 365.94 389.88 ;
   RECT 0.0 389.88 365.94 391.59 ;
   RECT 0.0 391.59 365.94 393.3 ;
   RECT 0.0 393.3 365.94 395.01 ;
   RECT 0.0 395.01 365.94 396.72 ;
   RECT 0.0 396.72 365.94 398.43 ;
   RECT 0.0 398.43 365.94 400.14 ;
   RECT 0.0 400.14 365.94 401.85 ;
   RECT 0.0 401.85 365.94 403.56 ;
   RECT 0.0 403.56 365.94 405.27 ;
   RECT 0.0 405.27 365.94 406.98 ;
   RECT 0.0 406.98 365.94 408.69 ;
   RECT 0.0 408.69 365.94 410.4 ;
   RECT 0.0 410.4 365.94 412.11 ;
   RECT 0.0 412.11 365.94 413.82 ;
   RECT 0.0 413.82 365.94 415.53 ;
   RECT 0.0 415.53 365.94 417.24 ;
   RECT 0.0 417.24 365.94 418.95 ;
   RECT 0.0 418.95 365.94 420.66 ;
   RECT 0.0 420.66 365.94 422.37 ;
   RECT 0.0 422.37 365.94 424.08 ;
   RECT 0.0 424.08 365.94 425.79 ;
   RECT 0.0 425.79 365.94 427.5 ;
   RECT 0.0 427.5 365.94 429.21 ;
   RECT 0.0 429.21 365.94 430.92 ;
   RECT 0.0 430.92 365.94 432.63 ;
   RECT 0.0 432.63 365.94 434.34 ;
   RECT 0.0 434.34 365.94 436.05 ;
   RECT 0.0 436.05 365.94 437.76 ;
   RECT 0.0 437.76 365.94 439.47 ;
   RECT 0.0 439.47 365.94 441.18 ;
   RECT 0.0 441.18 365.94 442.89 ;
   RECT 0.0 442.89 365.94 444.6 ;
   RECT 0.0 444.6 365.94 446.31 ;
   RECT 0.0 446.31 365.94 448.02 ;
   RECT 0.0 448.02 365.94 449.73 ;
   RECT 0.0 449.73 365.94 451.44 ;
   RECT 0.0 451.44 365.94 453.15 ;
   RECT 0.0 453.15 365.94 454.86 ;
   RECT 0.0 454.86 365.94 456.57 ;
   RECT 0.0 456.57 365.94 458.28 ;
   RECT 0.0 458.28 365.94 459.99 ;
   RECT 0.0 459.99 365.94 461.7 ;
   RECT 0.0 461.7 365.94 463.41 ;
   RECT 0.0 463.41 365.94 465.12 ;
   RECT 0.0 465.12 365.94 466.83 ;
   RECT 0.0 466.83 365.94 468.54 ;
   RECT 0.0 468.54 365.94 470.25 ;
   RECT 0.0 470.25 365.94 471.96 ;
   RECT 0.0 471.96 365.94 473.67 ;
   RECT 0.0 473.67 365.94 475.38 ;
  LAYER via1 ;
   RECT 0.0 0.0 365.94 1.71 ;
   RECT 0.0 1.71 365.94 3.42 ;
   RECT 0.0 3.42 365.94 5.13 ;
   RECT 0.0 5.13 365.94 6.84 ;
   RECT 0.0 6.84 365.94 8.55 ;
   RECT 0.0 8.55 365.94 10.26 ;
   RECT 0.0 10.26 365.94 11.97 ;
   RECT 0.0 11.97 365.94 13.68 ;
   RECT 0.0 13.68 365.94 15.39 ;
   RECT 0.0 15.39 365.94 17.1 ;
   RECT 0.0 17.1 365.94 18.81 ;
   RECT 0.0 18.81 365.94 20.52 ;
   RECT 0.0 20.52 365.94 22.23 ;
   RECT 0.0 22.23 365.94 23.94 ;
   RECT 0.0 23.94 365.94 25.65 ;
   RECT 0.0 25.65 365.94 27.36 ;
   RECT 0.0 27.36 365.94 29.07 ;
   RECT 0.0 29.07 365.94 30.78 ;
   RECT 0.0 30.78 365.94 32.49 ;
   RECT 0.0 32.49 365.94 34.2 ;
   RECT 0.0 34.2 365.94 35.91 ;
   RECT 0.0 35.91 365.94 37.62 ;
   RECT 0.0 37.62 365.94 39.33 ;
   RECT 0.0 39.33 365.94 41.04 ;
   RECT 0.0 41.04 365.94 42.75 ;
   RECT 0.0 42.75 365.94 44.46 ;
   RECT 0.0 44.46 365.94 46.17 ;
   RECT 0.0 46.17 365.94 47.88 ;
   RECT 0.0 47.88 365.94 49.59 ;
   RECT 0.0 49.59 365.94 51.3 ;
   RECT 0.0 51.3 365.94 53.01 ;
   RECT 0.0 53.01 365.94 54.72 ;
   RECT 0.0 54.72 365.94 56.43 ;
   RECT 0.0 56.43 365.94 58.14 ;
   RECT 0.0 58.14 365.94 59.85 ;
   RECT 0.0 59.85 365.94 61.56 ;
   RECT 0.0 61.56 365.94 63.27 ;
   RECT 0.0 63.27 365.94 64.98 ;
   RECT 0.0 64.98 365.94 66.69 ;
   RECT 0.0 66.69 365.94 68.4 ;
   RECT 0.0 68.4 365.94 70.11 ;
   RECT 0.0 70.11 365.94 71.82 ;
   RECT 0.0 71.82 365.94 73.53 ;
   RECT 0.0 73.53 365.94 75.24 ;
   RECT 0.0 75.24 365.94 76.95 ;
   RECT 0.0 76.95 365.94 78.66 ;
   RECT 0.0 78.66 365.94 80.37 ;
   RECT 0.0 80.37 365.94 82.08 ;
   RECT 0.0 82.08 365.94 83.79 ;
   RECT 0.0 83.79 365.94 85.5 ;
   RECT 0.0 85.5 365.94 87.21 ;
   RECT 0.0 87.21 365.94 88.92 ;
   RECT 0.0 88.92 365.94 90.63 ;
   RECT 0.0 90.63 365.94 92.34 ;
   RECT 0.0 92.34 365.94 94.05 ;
   RECT 0.0 94.05 365.94 95.76 ;
   RECT 0.0 95.76 365.94 97.47 ;
   RECT 0.0 97.47 365.94 99.18 ;
   RECT 0.0 99.18 365.94 100.89 ;
   RECT 0.0 100.89 365.94 102.6 ;
   RECT 0.0 102.6 365.94 104.31 ;
   RECT 0.0 104.31 365.94 106.02 ;
   RECT 0.0 106.02 365.94 107.73 ;
   RECT 0.0 107.73 365.94 109.44 ;
   RECT 0.0 109.44 365.94 111.15 ;
   RECT 0.0 111.15 365.94 112.86 ;
   RECT 0.0 112.86 365.94 114.57 ;
   RECT 0.0 114.57 365.94 116.28 ;
   RECT 0.0 116.28 365.94 117.99 ;
   RECT 0.0 117.99 365.94 119.7 ;
   RECT 0.0 119.7 365.94 121.41 ;
   RECT 0.0 121.41 365.94 123.12 ;
   RECT 0.0 123.12 365.94 124.83 ;
   RECT 0.0 124.83 365.94 126.54 ;
   RECT 0.0 126.54 365.94 128.25 ;
   RECT 0.0 128.25 365.94 129.96 ;
   RECT 0.0 129.96 365.94 131.67 ;
   RECT 0.0 131.67 365.94 133.38 ;
   RECT 0.0 133.38 365.94 135.09 ;
   RECT 0.0 135.09 365.94 136.8 ;
   RECT 0.0 136.8 365.94 138.51 ;
   RECT 0.0 138.51 365.94 140.22 ;
   RECT 0.0 140.22 365.94 141.93 ;
   RECT 0.0 141.93 365.94 143.64 ;
   RECT 0.0 143.64 365.94 145.35 ;
   RECT 0.0 145.35 365.94 147.06 ;
   RECT 0.0 147.06 365.94 148.77 ;
   RECT 0.0 148.77 365.94 150.48 ;
   RECT 0.0 150.48 365.94 152.19 ;
   RECT 0.0 152.19 365.94 153.9 ;
   RECT 0.0 153.9 365.94 155.61 ;
   RECT 0.0 155.61 365.94 157.32 ;
   RECT 0.0 157.32 365.94 159.03 ;
   RECT 0.0 159.03 365.94 160.74 ;
   RECT 0.0 160.74 365.94 162.45 ;
   RECT 0.0 162.45 365.94 164.16 ;
   RECT 0.0 164.16 365.94 165.87 ;
   RECT 0.0 165.87 365.94 167.58 ;
   RECT 0.0 167.58 365.94 169.29 ;
   RECT 0.0 169.29 365.94 171.0 ;
   RECT 0.0 171.0 365.94 172.71 ;
   RECT 0.0 172.71 365.94 174.42 ;
   RECT 0.0 174.42 365.94 176.13 ;
   RECT 0.0 176.13 365.94 177.84 ;
   RECT 0.0 177.84 365.94 179.55 ;
   RECT 0.0 179.55 365.94 181.26 ;
   RECT 0.0 181.26 365.94 182.97 ;
   RECT 0.0 182.97 365.94 184.68 ;
   RECT 0.0 184.68 365.94 186.39 ;
   RECT 0.0 186.39 365.94 188.1 ;
   RECT 0.0 188.1 365.94 189.81 ;
   RECT 0.0 189.81 365.94 191.52 ;
   RECT 0.0 191.52 365.94 193.23 ;
   RECT 0.0 193.23 365.94 194.94 ;
   RECT 0.0 194.94 365.94 196.65 ;
   RECT 0.0 196.65 365.94 198.36 ;
   RECT 0.0 198.36 365.94 200.07 ;
   RECT 0.0 200.07 365.94 201.78 ;
   RECT 0.0 201.78 365.94 203.49 ;
   RECT 0.0 203.49 365.94 205.2 ;
   RECT 0.0 205.2 365.94 206.91 ;
   RECT 0.0 206.91 365.94 208.62 ;
   RECT 0.0 208.62 365.94 210.33 ;
   RECT 0.0 210.33 365.94 212.04 ;
   RECT 0.0 212.04 365.94 213.75 ;
   RECT 0.0 213.75 365.94 215.46 ;
   RECT 0.0 215.46 365.94 217.17 ;
   RECT 0.0 217.17 365.94 218.88 ;
   RECT 0.0 218.88 365.94 220.59 ;
   RECT 0.0 220.59 365.94 222.3 ;
   RECT 0.0 222.3 365.94 224.01 ;
   RECT 0.0 224.01 365.94 225.72 ;
   RECT 0.0 225.72 365.94 227.43 ;
   RECT 0.0 227.43 365.94 229.14 ;
   RECT 0.0 229.14 365.94 230.85 ;
   RECT 0.0 230.85 389.12 232.56 ;
   RECT 0.0 232.56 389.12 234.27 ;
   RECT 0.0 234.27 389.12 235.98 ;
   RECT 0.0 235.98 389.12 237.69 ;
   RECT 0.0 237.69 389.12 239.4 ;
   RECT 0.0 239.4 389.12 241.11 ;
   RECT 0.0 241.11 389.12 242.82 ;
   RECT 0.0 242.82 389.12 244.53 ;
   RECT 0.0 244.53 389.12 246.24 ;
   RECT 0.0 246.24 389.12 247.95 ;
   RECT 0.0 247.95 389.12 249.66 ;
   RECT 0.0 249.66 389.12 251.37 ;
   RECT 0.0 251.37 389.12 253.08 ;
   RECT 0.0 253.08 389.12 254.79 ;
   RECT 0.0 254.79 389.12 256.5 ;
   RECT 0.0 256.5 389.12 258.21 ;
   RECT 0.0 258.21 389.12 259.92 ;
   RECT 0.0 259.92 365.94 261.63 ;
   RECT 0.0 261.63 365.94 263.34 ;
   RECT 0.0 263.34 365.94 265.05 ;
   RECT 0.0 265.05 365.94 266.76 ;
   RECT 0.0 266.76 365.94 268.47 ;
   RECT 0.0 268.47 365.94 270.18 ;
   RECT 0.0 270.18 365.94 271.89 ;
   RECT 0.0 271.89 365.94 273.6 ;
   RECT 0.0 273.6 365.94 275.31 ;
   RECT 0.0 275.31 365.94 277.02 ;
   RECT 0.0 277.02 365.94 278.73 ;
   RECT 0.0 278.73 365.94 280.44 ;
   RECT 0.0 280.44 365.94 282.15 ;
   RECT 0.0 282.15 365.94 283.86 ;
   RECT 0.0 283.86 365.94 285.57 ;
   RECT 0.0 285.57 365.94 287.28 ;
   RECT 0.0 287.28 365.94 288.99 ;
   RECT 0.0 288.99 365.94 290.7 ;
   RECT 0.0 290.7 365.94 292.41 ;
   RECT 0.0 292.41 365.94 294.12 ;
   RECT 0.0 294.12 365.94 295.83 ;
   RECT 0.0 295.83 365.94 297.54 ;
   RECT 0.0 297.54 365.94 299.25 ;
   RECT 0.0 299.25 365.94 300.96 ;
   RECT 0.0 300.96 365.94 302.67 ;
   RECT 0.0 302.67 365.94 304.38 ;
   RECT 0.0 304.38 365.94 306.09 ;
   RECT 0.0 306.09 365.94 307.8 ;
   RECT 0.0 307.8 365.94 309.51 ;
   RECT 0.0 309.51 365.94 311.22 ;
   RECT 0.0 311.22 365.94 312.93 ;
   RECT 0.0 312.93 365.94 314.64 ;
   RECT 0.0 314.64 365.94 316.35 ;
   RECT 0.0 316.35 365.94 318.06 ;
   RECT 0.0 318.06 365.94 319.77 ;
   RECT 0.0 319.77 365.94 321.48 ;
   RECT 0.0 321.48 365.94 323.19 ;
   RECT 0.0 323.19 365.94 324.9 ;
   RECT 0.0 324.9 365.94 326.61 ;
   RECT 0.0 326.61 365.94 328.32 ;
   RECT 0.0 328.32 365.94 330.03 ;
   RECT 0.0 330.03 365.94 331.74 ;
   RECT 0.0 331.74 365.94 333.45 ;
   RECT 0.0 333.45 365.94 335.16 ;
   RECT 0.0 335.16 365.94 336.87 ;
   RECT 0.0 336.87 365.94 338.58 ;
   RECT 0.0 338.58 365.94 340.29 ;
   RECT 0.0 340.29 365.94 342.0 ;
   RECT 0.0 342.0 365.94 343.71 ;
   RECT 0.0 343.71 365.94 345.42 ;
   RECT 0.0 345.42 365.94 347.13 ;
   RECT 0.0 347.13 365.94 348.84 ;
   RECT 0.0 348.84 365.94 350.55 ;
   RECT 0.0 350.55 365.94 352.26 ;
   RECT 0.0 352.26 365.94 353.97 ;
   RECT 0.0 353.97 365.94 355.68 ;
   RECT 0.0 355.68 365.94 357.39 ;
   RECT 0.0 357.39 365.94 359.1 ;
   RECT 0.0 359.1 365.94 360.81 ;
   RECT 0.0 360.81 365.94 362.52 ;
   RECT 0.0 362.52 365.94 364.23 ;
   RECT 0.0 364.23 365.94 365.94 ;
   RECT 0.0 365.94 365.94 367.65 ;
   RECT 0.0 367.65 365.94 369.36 ;
   RECT 0.0 369.36 365.94 371.07 ;
   RECT 0.0 371.07 365.94 372.78 ;
   RECT 0.0 372.78 365.94 374.49 ;
   RECT 0.0 374.49 365.94 376.2 ;
   RECT 0.0 376.2 365.94 377.91 ;
   RECT 0.0 377.91 365.94 379.62 ;
   RECT 0.0 379.62 365.94 381.33 ;
   RECT 0.0 381.33 365.94 383.04 ;
   RECT 0.0 383.04 365.94 384.75 ;
   RECT 0.0 384.75 365.94 386.46 ;
   RECT 0.0 386.46 365.94 388.17 ;
   RECT 0.0 388.17 365.94 389.88 ;
   RECT 0.0 389.88 365.94 391.59 ;
   RECT 0.0 391.59 365.94 393.3 ;
   RECT 0.0 393.3 365.94 395.01 ;
   RECT 0.0 395.01 365.94 396.72 ;
   RECT 0.0 396.72 365.94 398.43 ;
   RECT 0.0 398.43 365.94 400.14 ;
   RECT 0.0 400.14 365.94 401.85 ;
   RECT 0.0 401.85 365.94 403.56 ;
   RECT 0.0 403.56 365.94 405.27 ;
   RECT 0.0 405.27 365.94 406.98 ;
   RECT 0.0 406.98 365.94 408.69 ;
   RECT 0.0 408.69 365.94 410.4 ;
   RECT 0.0 410.4 365.94 412.11 ;
   RECT 0.0 412.11 365.94 413.82 ;
   RECT 0.0 413.82 365.94 415.53 ;
   RECT 0.0 415.53 365.94 417.24 ;
   RECT 0.0 417.24 365.94 418.95 ;
   RECT 0.0 418.95 365.94 420.66 ;
   RECT 0.0 420.66 365.94 422.37 ;
   RECT 0.0 422.37 365.94 424.08 ;
   RECT 0.0 424.08 365.94 425.79 ;
   RECT 0.0 425.79 365.94 427.5 ;
   RECT 0.0 427.5 365.94 429.21 ;
   RECT 0.0 429.21 365.94 430.92 ;
   RECT 0.0 430.92 365.94 432.63 ;
   RECT 0.0 432.63 365.94 434.34 ;
   RECT 0.0 434.34 365.94 436.05 ;
   RECT 0.0 436.05 365.94 437.76 ;
   RECT 0.0 437.76 365.94 439.47 ;
   RECT 0.0 439.47 365.94 441.18 ;
   RECT 0.0 441.18 365.94 442.89 ;
   RECT 0.0 442.89 365.94 444.6 ;
   RECT 0.0 444.6 365.94 446.31 ;
   RECT 0.0 446.31 365.94 448.02 ;
   RECT 0.0 448.02 365.94 449.73 ;
   RECT 0.0 449.73 365.94 451.44 ;
   RECT 0.0 451.44 365.94 453.15 ;
   RECT 0.0 453.15 365.94 454.86 ;
   RECT 0.0 454.86 365.94 456.57 ;
   RECT 0.0 456.57 365.94 458.28 ;
   RECT 0.0 458.28 365.94 459.99 ;
   RECT 0.0 459.99 365.94 461.7 ;
   RECT 0.0 461.7 365.94 463.41 ;
   RECT 0.0 463.41 365.94 465.12 ;
   RECT 0.0 465.12 365.94 466.83 ;
   RECT 0.0 466.83 365.94 468.54 ;
   RECT 0.0 468.54 365.94 470.25 ;
   RECT 0.0 470.25 365.94 471.96 ;
   RECT 0.0 471.96 365.94 473.67 ;
   RECT 0.0 473.67 365.94 475.38 ;
  LAYER metal2 ;
   RECT 0.0 0.0 365.94 1.71 ;
   RECT 0.0 1.71 365.94 3.42 ;
   RECT 0.0 3.42 365.94 5.13 ;
   RECT 0.0 5.13 365.94 6.84 ;
   RECT 0.0 6.84 365.94 8.55 ;
   RECT 0.0 8.55 365.94 10.26 ;
   RECT 0.0 10.26 365.94 11.97 ;
   RECT 0.0 11.97 365.94 13.68 ;
   RECT 0.0 13.68 365.94 15.39 ;
   RECT 0.0 15.39 365.94 17.1 ;
   RECT 0.0 17.1 365.94 18.81 ;
   RECT 0.0 18.81 365.94 20.52 ;
   RECT 0.0 20.52 365.94 22.23 ;
   RECT 0.0 22.23 365.94 23.94 ;
   RECT 0.0 23.94 365.94 25.65 ;
   RECT 0.0 25.65 365.94 27.36 ;
   RECT 0.0 27.36 365.94 29.07 ;
   RECT 0.0 29.07 365.94 30.78 ;
   RECT 0.0 30.78 365.94 32.49 ;
   RECT 0.0 32.49 365.94 34.2 ;
   RECT 0.0 34.2 365.94 35.91 ;
   RECT 0.0 35.91 365.94 37.62 ;
   RECT 0.0 37.62 365.94 39.33 ;
   RECT 0.0 39.33 365.94 41.04 ;
   RECT 0.0 41.04 365.94 42.75 ;
   RECT 0.0 42.75 365.94 44.46 ;
   RECT 0.0 44.46 365.94 46.17 ;
   RECT 0.0 46.17 365.94 47.88 ;
   RECT 0.0 47.88 365.94 49.59 ;
   RECT 0.0 49.59 365.94 51.3 ;
   RECT 0.0 51.3 365.94 53.01 ;
   RECT 0.0 53.01 365.94 54.72 ;
   RECT 0.0 54.72 365.94 56.43 ;
   RECT 0.0 56.43 365.94 58.14 ;
   RECT 0.0 58.14 365.94 59.85 ;
   RECT 0.0 59.85 365.94 61.56 ;
   RECT 0.0 61.56 365.94 63.27 ;
   RECT 0.0 63.27 365.94 64.98 ;
   RECT 0.0 64.98 365.94 66.69 ;
   RECT 0.0 66.69 365.94 68.4 ;
   RECT 0.0 68.4 365.94 70.11 ;
   RECT 0.0 70.11 365.94 71.82 ;
   RECT 0.0 71.82 365.94 73.53 ;
   RECT 0.0 73.53 365.94 75.24 ;
   RECT 0.0 75.24 365.94 76.95 ;
   RECT 0.0 76.95 365.94 78.66 ;
   RECT 0.0 78.66 365.94 80.37 ;
   RECT 0.0 80.37 365.94 82.08 ;
   RECT 0.0 82.08 365.94 83.79 ;
   RECT 0.0 83.79 365.94 85.5 ;
   RECT 0.0 85.5 365.94 87.21 ;
   RECT 0.0 87.21 365.94 88.92 ;
   RECT 0.0 88.92 365.94 90.63 ;
   RECT 0.0 90.63 365.94 92.34 ;
   RECT 0.0 92.34 365.94 94.05 ;
   RECT 0.0 94.05 365.94 95.76 ;
   RECT 0.0 95.76 365.94 97.47 ;
   RECT 0.0 97.47 365.94 99.18 ;
   RECT 0.0 99.18 365.94 100.89 ;
   RECT 0.0 100.89 365.94 102.6 ;
   RECT 0.0 102.6 365.94 104.31 ;
   RECT 0.0 104.31 365.94 106.02 ;
   RECT 0.0 106.02 365.94 107.73 ;
   RECT 0.0 107.73 365.94 109.44 ;
   RECT 0.0 109.44 365.94 111.15 ;
   RECT 0.0 111.15 365.94 112.86 ;
   RECT 0.0 112.86 365.94 114.57 ;
   RECT 0.0 114.57 365.94 116.28 ;
   RECT 0.0 116.28 365.94 117.99 ;
   RECT 0.0 117.99 365.94 119.7 ;
   RECT 0.0 119.7 365.94 121.41 ;
   RECT 0.0 121.41 365.94 123.12 ;
   RECT 0.0 123.12 365.94 124.83 ;
   RECT 0.0 124.83 365.94 126.54 ;
   RECT 0.0 126.54 365.94 128.25 ;
   RECT 0.0 128.25 365.94 129.96 ;
   RECT 0.0 129.96 365.94 131.67 ;
   RECT 0.0 131.67 365.94 133.38 ;
   RECT 0.0 133.38 365.94 135.09 ;
   RECT 0.0 135.09 365.94 136.8 ;
   RECT 0.0 136.8 365.94 138.51 ;
   RECT 0.0 138.51 365.94 140.22 ;
   RECT 0.0 140.22 365.94 141.93 ;
   RECT 0.0 141.93 365.94 143.64 ;
   RECT 0.0 143.64 365.94 145.35 ;
   RECT 0.0 145.35 365.94 147.06 ;
   RECT 0.0 147.06 365.94 148.77 ;
   RECT 0.0 148.77 365.94 150.48 ;
   RECT 0.0 150.48 365.94 152.19 ;
   RECT 0.0 152.19 365.94 153.9 ;
   RECT 0.0 153.9 365.94 155.61 ;
   RECT 0.0 155.61 365.94 157.32 ;
   RECT 0.0 157.32 365.94 159.03 ;
   RECT 0.0 159.03 365.94 160.74 ;
   RECT 0.0 160.74 365.94 162.45 ;
   RECT 0.0 162.45 365.94 164.16 ;
   RECT 0.0 164.16 365.94 165.87 ;
   RECT 0.0 165.87 365.94 167.58 ;
   RECT 0.0 167.58 365.94 169.29 ;
   RECT 0.0 169.29 365.94 171.0 ;
   RECT 0.0 171.0 365.94 172.71 ;
   RECT 0.0 172.71 365.94 174.42 ;
   RECT 0.0 174.42 365.94 176.13 ;
   RECT 0.0 176.13 365.94 177.84 ;
   RECT 0.0 177.84 365.94 179.55 ;
   RECT 0.0 179.55 365.94 181.26 ;
   RECT 0.0 181.26 365.94 182.97 ;
   RECT 0.0 182.97 365.94 184.68 ;
   RECT 0.0 184.68 365.94 186.39 ;
   RECT 0.0 186.39 365.94 188.1 ;
   RECT 0.0 188.1 365.94 189.81 ;
   RECT 0.0 189.81 365.94 191.52 ;
   RECT 0.0 191.52 365.94 193.23 ;
   RECT 0.0 193.23 365.94 194.94 ;
   RECT 0.0 194.94 365.94 196.65 ;
   RECT 0.0 196.65 365.94 198.36 ;
   RECT 0.0 198.36 365.94 200.07 ;
   RECT 0.0 200.07 365.94 201.78 ;
   RECT 0.0 201.78 365.94 203.49 ;
   RECT 0.0 203.49 365.94 205.2 ;
   RECT 0.0 205.2 365.94 206.91 ;
   RECT 0.0 206.91 365.94 208.62 ;
   RECT 0.0 208.62 365.94 210.33 ;
   RECT 0.0 210.33 365.94 212.04 ;
   RECT 0.0 212.04 365.94 213.75 ;
   RECT 0.0 213.75 365.94 215.46 ;
   RECT 0.0 215.46 365.94 217.17 ;
   RECT 0.0 217.17 365.94 218.88 ;
   RECT 0.0 218.88 365.94 220.59 ;
   RECT 0.0 220.59 365.94 222.3 ;
   RECT 0.0 222.3 365.94 224.01 ;
   RECT 0.0 224.01 365.94 225.72 ;
   RECT 0.0 225.72 365.94 227.43 ;
   RECT 0.0 227.43 365.94 229.14 ;
   RECT 0.0 229.14 365.94 230.85 ;
   RECT 0.0 230.85 389.12 232.56 ;
   RECT 0.0 232.56 389.12 234.27 ;
   RECT 0.0 234.27 389.12 235.98 ;
   RECT 0.0 235.98 389.12 237.69 ;
   RECT 0.0 237.69 389.12 239.4 ;
   RECT 0.0 239.4 389.12 241.11 ;
   RECT 0.0 241.11 389.12 242.82 ;
   RECT 0.0 242.82 389.12 244.53 ;
   RECT 0.0 244.53 389.12 246.24 ;
   RECT 0.0 246.24 389.12 247.95 ;
   RECT 0.0 247.95 389.12 249.66 ;
   RECT 0.0 249.66 389.12 251.37 ;
   RECT 0.0 251.37 389.12 253.08 ;
   RECT 0.0 253.08 389.12 254.79 ;
   RECT 0.0 254.79 389.12 256.5 ;
   RECT 0.0 256.5 389.12 258.21 ;
   RECT 0.0 258.21 389.12 259.92 ;
   RECT 0.0 259.92 365.94 261.63 ;
   RECT 0.0 261.63 365.94 263.34 ;
   RECT 0.0 263.34 365.94 265.05 ;
   RECT 0.0 265.05 365.94 266.76 ;
   RECT 0.0 266.76 365.94 268.47 ;
   RECT 0.0 268.47 365.94 270.18 ;
   RECT 0.0 270.18 365.94 271.89 ;
   RECT 0.0 271.89 365.94 273.6 ;
   RECT 0.0 273.6 365.94 275.31 ;
   RECT 0.0 275.31 365.94 277.02 ;
   RECT 0.0 277.02 365.94 278.73 ;
   RECT 0.0 278.73 365.94 280.44 ;
   RECT 0.0 280.44 365.94 282.15 ;
   RECT 0.0 282.15 365.94 283.86 ;
   RECT 0.0 283.86 365.94 285.57 ;
   RECT 0.0 285.57 365.94 287.28 ;
   RECT 0.0 287.28 365.94 288.99 ;
   RECT 0.0 288.99 365.94 290.7 ;
   RECT 0.0 290.7 365.94 292.41 ;
   RECT 0.0 292.41 365.94 294.12 ;
   RECT 0.0 294.12 365.94 295.83 ;
   RECT 0.0 295.83 365.94 297.54 ;
   RECT 0.0 297.54 365.94 299.25 ;
   RECT 0.0 299.25 365.94 300.96 ;
   RECT 0.0 300.96 365.94 302.67 ;
   RECT 0.0 302.67 365.94 304.38 ;
   RECT 0.0 304.38 365.94 306.09 ;
   RECT 0.0 306.09 365.94 307.8 ;
   RECT 0.0 307.8 365.94 309.51 ;
   RECT 0.0 309.51 365.94 311.22 ;
   RECT 0.0 311.22 365.94 312.93 ;
   RECT 0.0 312.93 365.94 314.64 ;
   RECT 0.0 314.64 365.94 316.35 ;
   RECT 0.0 316.35 365.94 318.06 ;
   RECT 0.0 318.06 365.94 319.77 ;
   RECT 0.0 319.77 365.94 321.48 ;
   RECT 0.0 321.48 365.94 323.19 ;
   RECT 0.0 323.19 365.94 324.9 ;
   RECT 0.0 324.9 365.94 326.61 ;
   RECT 0.0 326.61 365.94 328.32 ;
   RECT 0.0 328.32 365.94 330.03 ;
   RECT 0.0 330.03 365.94 331.74 ;
   RECT 0.0 331.74 365.94 333.45 ;
   RECT 0.0 333.45 365.94 335.16 ;
   RECT 0.0 335.16 365.94 336.87 ;
   RECT 0.0 336.87 365.94 338.58 ;
   RECT 0.0 338.58 365.94 340.29 ;
   RECT 0.0 340.29 365.94 342.0 ;
   RECT 0.0 342.0 365.94 343.71 ;
   RECT 0.0 343.71 365.94 345.42 ;
   RECT 0.0 345.42 365.94 347.13 ;
   RECT 0.0 347.13 365.94 348.84 ;
   RECT 0.0 348.84 365.94 350.55 ;
   RECT 0.0 350.55 365.94 352.26 ;
   RECT 0.0 352.26 365.94 353.97 ;
   RECT 0.0 353.97 365.94 355.68 ;
   RECT 0.0 355.68 365.94 357.39 ;
   RECT 0.0 357.39 365.94 359.1 ;
   RECT 0.0 359.1 365.94 360.81 ;
   RECT 0.0 360.81 365.94 362.52 ;
   RECT 0.0 362.52 365.94 364.23 ;
   RECT 0.0 364.23 365.94 365.94 ;
   RECT 0.0 365.94 365.94 367.65 ;
   RECT 0.0 367.65 365.94 369.36 ;
   RECT 0.0 369.36 365.94 371.07 ;
   RECT 0.0 371.07 365.94 372.78 ;
   RECT 0.0 372.78 365.94 374.49 ;
   RECT 0.0 374.49 365.94 376.2 ;
   RECT 0.0 376.2 365.94 377.91 ;
   RECT 0.0 377.91 365.94 379.62 ;
   RECT 0.0 379.62 365.94 381.33 ;
   RECT 0.0 381.33 365.94 383.04 ;
   RECT 0.0 383.04 365.94 384.75 ;
   RECT 0.0 384.75 365.94 386.46 ;
   RECT 0.0 386.46 365.94 388.17 ;
   RECT 0.0 388.17 365.94 389.88 ;
   RECT 0.0 389.88 365.94 391.59 ;
   RECT 0.0 391.59 365.94 393.3 ;
   RECT 0.0 393.3 365.94 395.01 ;
   RECT 0.0 395.01 365.94 396.72 ;
   RECT 0.0 396.72 365.94 398.43 ;
   RECT 0.0 398.43 365.94 400.14 ;
   RECT 0.0 400.14 365.94 401.85 ;
   RECT 0.0 401.85 365.94 403.56 ;
   RECT 0.0 403.56 365.94 405.27 ;
   RECT 0.0 405.27 365.94 406.98 ;
   RECT 0.0 406.98 365.94 408.69 ;
   RECT 0.0 408.69 365.94 410.4 ;
   RECT 0.0 410.4 365.94 412.11 ;
   RECT 0.0 412.11 365.94 413.82 ;
   RECT 0.0 413.82 365.94 415.53 ;
   RECT 0.0 415.53 365.94 417.24 ;
   RECT 0.0 417.24 365.94 418.95 ;
   RECT 0.0 418.95 365.94 420.66 ;
   RECT 0.0 420.66 365.94 422.37 ;
   RECT 0.0 422.37 365.94 424.08 ;
   RECT 0.0 424.08 365.94 425.79 ;
   RECT 0.0 425.79 365.94 427.5 ;
   RECT 0.0 427.5 365.94 429.21 ;
   RECT 0.0 429.21 365.94 430.92 ;
   RECT 0.0 430.92 365.94 432.63 ;
   RECT 0.0 432.63 365.94 434.34 ;
   RECT 0.0 434.34 365.94 436.05 ;
   RECT 0.0 436.05 365.94 437.76 ;
   RECT 0.0 437.76 365.94 439.47 ;
   RECT 0.0 439.47 365.94 441.18 ;
   RECT 0.0 441.18 365.94 442.89 ;
   RECT 0.0 442.89 365.94 444.6 ;
   RECT 0.0 444.6 365.94 446.31 ;
   RECT 0.0 446.31 365.94 448.02 ;
   RECT 0.0 448.02 365.94 449.73 ;
   RECT 0.0 449.73 365.94 451.44 ;
   RECT 0.0 451.44 365.94 453.15 ;
   RECT 0.0 453.15 365.94 454.86 ;
   RECT 0.0 454.86 365.94 456.57 ;
   RECT 0.0 456.57 365.94 458.28 ;
   RECT 0.0 458.28 365.94 459.99 ;
   RECT 0.0 459.99 365.94 461.7 ;
   RECT 0.0 461.7 365.94 463.41 ;
   RECT 0.0 463.41 365.94 465.12 ;
   RECT 0.0 465.12 365.94 466.83 ;
   RECT 0.0 466.83 365.94 468.54 ;
   RECT 0.0 468.54 365.94 470.25 ;
   RECT 0.0 470.25 365.94 471.96 ;
   RECT 0.0 471.96 365.94 473.67 ;
   RECT 0.0 473.67 365.94 475.38 ;
  LAYER via2 ;
   RECT 0.0 0.0 365.94 1.71 ;
   RECT 0.0 1.71 365.94 3.42 ;
   RECT 0.0 3.42 365.94 5.13 ;
   RECT 0.0 5.13 365.94 6.84 ;
   RECT 0.0 6.84 365.94 8.55 ;
   RECT 0.0 8.55 365.94 10.26 ;
   RECT 0.0 10.26 365.94 11.97 ;
   RECT 0.0 11.97 365.94 13.68 ;
   RECT 0.0 13.68 365.94 15.39 ;
   RECT 0.0 15.39 365.94 17.1 ;
   RECT 0.0 17.1 365.94 18.81 ;
   RECT 0.0 18.81 365.94 20.52 ;
   RECT 0.0 20.52 365.94 22.23 ;
   RECT 0.0 22.23 365.94 23.94 ;
   RECT 0.0 23.94 365.94 25.65 ;
   RECT 0.0 25.65 365.94 27.36 ;
   RECT 0.0 27.36 365.94 29.07 ;
   RECT 0.0 29.07 365.94 30.78 ;
   RECT 0.0 30.78 365.94 32.49 ;
   RECT 0.0 32.49 365.94 34.2 ;
   RECT 0.0 34.2 365.94 35.91 ;
   RECT 0.0 35.91 365.94 37.62 ;
   RECT 0.0 37.62 365.94 39.33 ;
   RECT 0.0 39.33 365.94 41.04 ;
   RECT 0.0 41.04 365.94 42.75 ;
   RECT 0.0 42.75 365.94 44.46 ;
   RECT 0.0 44.46 365.94 46.17 ;
   RECT 0.0 46.17 365.94 47.88 ;
   RECT 0.0 47.88 365.94 49.59 ;
   RECT 0.0 49.59 365.94 51.3 ;
   RECT 0.0 51.3 365.94 53.01 ;
   RECT 0.0 53.01 365.94 54.72 ;
   RECT 0.0 54.72 365.94 56.43 ;
   RECT 0.0 56.43 365.94 58.14 ;
   RECT 0.0 58.14 365.94 59.85 ;
   RECT 0.0 59.85 365.94 61.56 ;
   RECT 0.0 61.56 365.94 63.27 ;
   RECT 0.0 63.27 365.94 64.98 ;
   RECT 0.0 64.98 365.94 66.69 ;
   RECT 0.0 66.69 365.94 68.4 ;
   RECT 0.0 68.4 365.94 70.11 ;
   RECT 0.0 70.11 365.94 71.82 ;
   RECT 0.0 71.82 365.94 73.53 ;
   RECT 0.0 73.53 365.94 75.24 ;
   RECT 0.0 75.24 365.94 76.95 ;
   RECT 0.0 76.95 365.94 78.66 ;
   RECT 0.0 78.66 365.94 80.37 ;
   RECT 0.0 80.37 365.94 82.08 ;
   RECT 0.0 82.08 365.94 83.79 ;
   RECT 0.0 83.79 365.94 85.5 ;
   RECT 0.0 85.5 365.94 87.21 ;
   RECT 0.0 87.21 365.94 88.92 ;
   RECT 0.0 88.92 365.94 90.63 ;
   RECT 0.0 90.63 365.94 92.34 ;
   RECT 0.0 92.34 365.94 94.05 ;
   RECT 0.0 94.05 365.94 95.76 ;
   RECT 0.0 95.76 365.94 97.47 ;
   RECT 0.0 97.47 365.94 99.18 ;
   RECT 0.0 99.18 365.94 100.89 ;
   RECT 0.0 100.89 365.94 102.6 ;
   RECT 0.0 102.6 365.94 104.31 ;
   RECT 0.0 104.31 365.94 106.02 ;
   RECT 0.0 106.02 365.94 107.73 ;
   RECT 0.0 107.73 365.94 109.44 ;
   RECT 0.0 109.44 365.94 111.15 ;
   RECT 0.0 111.15 365.94 112.86 ;
   RECT 0.0 112.86 365.94 114.57 ;
   RECT 0.0 114.57 365.94 116.28 ;
   RECT 0.0 116.28 365.94 117.99 ;
   RECT 0.0 117.99 365.94 119.7 ;
   RECT 0.0 119.7 365.94 121.41 ;
   RECT 0.0 121.41 365.94 123.12 ;
   RECT 0.0 123.12 365.94 124.83 ;
   RECT 0.0 124.83 365.94 126.54 ;
   RECT 0.0 126.54 365.94 128.25 ;
   RECT 0.0 128.25 365.94 129.96 ;
   RECT 0.0 129.96 365.94 131.67 ;
   RECT 0.0 131.67 365.94 133.38 ;
   RECT 0.0 133.38 365.94 135.09 ;
   RECT 0.0 135.09 365.94 136.8 ;
   RECT 0.0 136.8 365.94 138.51 ;
   RECT 0.0 138.51 365.94 140.22 ;
   RECT 0.0 140.22 365.94 141.93 ;
   RECT 0.0 141.93 365.94 143.64 ;
   RECT 0.0 143.64 365.94 145.35 ;
   RECT 0.0 145.35 365.94 147.06 ;
   RECT 0.0 147.06 365.94 148.77 ;
   RECT 0.0 148.77 365.94 150.48 ;
   RECT 0.0 150.48 365.94 152.19 ;
   RECT 0.0 152.19 365.94 153.9 ;
   RECT 0.0 153.9 365.94 155.61 ;
   RECT 0.0 155.61 365.94 157.32 ;
   RECT 0.0 157.32 365.94 159.03 ;
   RECT 0.0 159.03 365.94 160.74 ;
   RECT 0.0 160.74 365.94 162.45 ;
   RECT 0.0 162.45 365.94 164.16 ;
   RECT 0.0 164.16 365.94 165.87 ;
   RECT 0.0 165.87 365.94 167.58 ;
   RECT 0.0 167.58 365.94 169.29 ;
   RECT 0.0 169.29 365.94 171.0 ;
   RECT 0.0 171.0 365.94 172.71 ;
   RECT 0.0 172.71 365.94 174.42 ;
   RECT 0.0 174.42 365.94 176.13 ;
   RECT 0.0 176.13 365.94 177.84 ;
   RECT 0.0 177.84 365.94 179.55 ;
   RECT 0.0 179.55 365.94 181.26 ;
   RECT 0.0 181.26 365.94 182.97 ;
   RECT 0.0 182.97 365.94 184.68 ;
   RECT 0.0 184.68 365.94 186.39 ;
   RECT 0.0 186.39 365.94 188.1 ;
   RECT 0.0 188.1 365.94 189.81 ;
   RECT 0.0 189.81 365.94 191.52 ;
   RECT 0.0 191.52 365.94 193.23 ;
   RECT 0.0 193.23 365.94 194.94 ;
   RECT 0.0 194.94 365.94 196.65 ;
   RECT 0.0 196.65 365.94 198.36 ;
   RECT 0.0 198.36 365.94 200.07 ;
   RECT 0.0 200.07 365.94 201.78 ;
   RECT 0.0 201.78 365.94 203.49 ;
   RECT 0.0 203.49 365.94 205.2 ;
   RECT 0.0 205.2 365.94 206.91 ;
   RECT 0.0 206.91 365.94 208.62 ;
   RECT 0.0 208.62 365.94 210.33 ;
   RECT 0.0 210.33 365.94 212.04 ;
   RECT 0.0 212.04 365.94 213.75 ;
   RECT 0.0 213.75 365.94 215.46 ;
   RECT 0.0 215.46 365.94 217.17 ;
   RECT 0.0 217.17 365.94 218.88 ;
   RECT 0.0 218.88 365.94 220.59 ;
   RECT 0.0 220.59 365.94 222.3 ;
   RECT 0.0 222.3 365.94 224.01 ;
   RECT 0.0 224.01 365.94 225.72 ;
   RECT 0.0 225.72 365.94 227.43 ;
   RECT 0.0 227.43 365.94 229.14 ;
   RECT 0.0 229.14 365.94 230.85 ;
   RECT 0.0 230.85 389.12 232.56 ;
   RECT 0.0 232.56 389.12 234.27 ;
   RECT 0.0 234.27 389.12 235.98 ;
   RECT 0.0 235.98 389.12 237.69 ;
   RECT 0.0 237.69 389.12 239.4 ;
   RECT 0.0 239.4 389.12 241.11 ;
   RECT 0.0 241.11 389.12 242.82 ;
   RECT 0.0 242.82 389.12 244.53 ;
   RECT 0.0 244.53 389.12 246.24 ;
   RECT 0.0 246.24 389.12 247.95 ;
   RECT 0.0 247.95 389.12 249.66 ;
   RECT 0.0 249.66 389.12 251.37 ;
   RECT 0.0 251.37 389.12 253.08 ;
   RECT 0.0 253.08 389.12 254.79 ;
   RECT 0.0 254.79 389.12 256.5 ;
   RECT 0.0 256.5 389.12 258.21 ;
   RECT 0.0 258.21 389.12 259.92 ;
   RECT 0.0 259.92 365.94 261.63 ;
   RECT 0.0 261.63 365.94 263.34 ;
   RECT 0.0 263.34 365.94 265.05 ;
   RECT 0.0 265.05 365.94 266.76 ;
   RECT 0.0 266.76 365.94 268.47 ;
   RECT 0.0 268.47 365.94 270.18 ;
   RECT 0.0 270.18 365.94 271.89 ;
   RECT 0.0 271.89 365.94 273.6 ;
   RECT 0.0 273.6 365.94 275.31 ;
   RECT 0.0 275.31 365.94 277.02 ;
   RECT 0.0 277.02 365.94 278.73 ;
   RECT 0.0 278.73 365.94 280.44 ;
   RECT 0.0 280.44 365.94 282.15 ;
   RECT 0.0 282.15 365.94 283.86 ;
   RECT 0.0 283.86 365.94 285.57 ;
   RECT 0.0 285.57 365.94 287.28 ;
   RECT 0.0 287.28 365.94 288.99 ;
   RECT 0.0 288.99 365.94 290.7 ;
   RECT 0.0 290.7 365.94 292.41 ;
   RECT 0.0 292.41 365.94 294.12 ;
   RECT 0.0 294.12 365.94 295.83 ;
   RECT 0.0 295.83 365.94 297.54 ;
   RECT 0.0 297.54 365.94 299.25 ;
   RECT 0.0 299.25 365.94 300.96 ;
   RECT 0.0 300.96 365.94 302.67 ;
   RECT 0.0 302.67 365.94 304.38 ;
   RECT 0.0 304.38 365.94 306.09 ;
   RECT 0.0 306.09 365.94 307.8 ;
   RECT 0.0 307.8 365.94 309.51 ;
   RECT 0.0 309.51 365.94 311.22 ;
   RECT 0.0 311.22 365.94 312.93 ;
   RECT 0.0 312.93 365.94 314.64 ;
   RECT 0.0 314.64 365.94 316.35 ;
   RECT 0.0 316.35 365.94 318.06 ;
   RECT 0.0 318.06 365.94 319.77 ;
   RECT 0.0 319.77 365.94 321.48 ;
   RECT 0.0 321.48 365.94 323.19 ;
   RECT 0.0 323.19 365.94 324.9 ;
   RECT 0.0 324.9 365.94 326.61 ;
   RECT 0.0 326.61 365.94 328.32 ;
   RECT 0.0 328.32 365.94 330.03 ;
   RECT 0.0 330.03 365.94 331.74 ;
   RECT 0.0 331.74 365.94 333.45 ;
   RECT 0.0 333.45 365.94 335.16 ;
   RECT 0.0 335.16 365.94 336.87 ;
   RECT 0.0 336.87 365.94 338.58 ;
   RECT 0.0 338.58 365.94 340.29 ;
   RECT 0.0 340.29 365.94 342.0 ;
   RECT 0.0 342.0 365.94 343.71 ;
   RECT 0.0 343.71 365.94 345.42 ;
   RECT 0.0 345.42 365.94 347.13 ;
   RECT 0.0 347.13 365.94 348.84 ;
   RECT 0.0 348.84 365.94 350.55 ;
   RECT 0.0 350.55 365.94 352.26 ;
   RECT 0.0 352.26 365.94 353.97 ;
   RECT 0.0 353.97 365.94 355.68 ;
   RECT 0.0 355.68 365.94 357.39 ;
   RECT 0.0 357.39 365.94 359.1 ;
   RECT 0.0 359.1 365.94 360.81 ;
   RECT 0.0 360.81 365.94 362.52 ;
   RECT 0.0 362.52 365.94 364.23 ;
   RECT 0.0 364.23 365.94 365.94 ;
   RECT 0.0 365.94 365.94 367.65 ;
   RECT 0.0 367.65 365.94 369.36 ;
   RECT 0.0 369.36 365.94 371.07 ;
   RECT 0.0 371.07 365.94 372.78 ;
   RECT 0.0 372.78 365.94 374.49 ;
   RECT 0.0 374.49 365.94 376.2 ;
   RECT 0.0 376.2 365.94 377.91 ;
   RECT 0.0 377.91 365.94 379.62 ;
   RECT 0.0 379.62 365.94 381.33 ;
   RECT 0.0 381.33 365.94 383.04 ;
   RECT 0.0 383.04 365.94 384.75 ;
   RECT 0.0 384.75 365.94 386.46 ;
   RECT 0.0 386.46 365.94 388.17 ;
   RECT 0.0 388.17 365.94 389.88 ;
   RECT 0.0 389.88 365.94 391.59 ;
   RECT 0.0 391.59 365.94 393.3 ;
   RECT 0.0 393.3 365.94 395.01 ;
   RECT 0.0 395.01 365.94 396.72 ;
   RECT 0.0 396.72 365.94 398.43 ;
   RECT 0.0 398.43 365.94 400.14 ;
   RECT 0.0 400.14 365.94 401.85 ;
   RECT 0.0 401.85 365.94 403.56 ;
   RECT 0.0 403.56 365.94 405.27 ;
   RECT 0.0 405.27 365.94 406.98 ;
   RECT 0.0 406.98 365.94 408.69 ;
   RECT 0.0 408.69 365.94 410.4 ;
   RECT 0.0 410.4 365.94 412.11 ;
   RECT 0.0 412.11 365.94 413.82 ;
   RECT 0.0 413.82 365.94 415.53 ;
   RECT 0.0 415.53 365.94 417.24 ;
   RECT 0.0 417.24 365.94 418.95 ;
   RECT 0.0 418.95 365.94 420.66 ;
   RECT 0.0 420.66 365.94 422.37 ;
   RECT 0.0 422.37 365.94 424.08 ;
   RECT 0.0 424.08 365.94 425.79 ;
   RECT 0.0 425.79 365.94 427.5 ;
   RECT 0.0 427.5 365.94 429.21 ;
   RECT 0.0 429.21 365.94 430.92 ;
   RECT 0.0 430.92 365.94 432.63 ;
   RECT 0.0 432.63 365.94 434.34 ;
   RECT 0.0 434.34 365.94 436.05 ;
   RECT 0.0 436.05 365.94 437.76 ;
   RECT 0.0 437.76 365.94 439.47 ;
   RECT 0.0 439.47 365.94 441.18 ;
   RECT 0.0 441.18 365.94 442.89 ;
   RECT 0.0 442.89 365.94 444.6 ;
   RECT 0.0 444.6 365.94 446.31 ;
   RECT 0.0 446.31 365.94 448.02 ;
   RECT 0.0 448.02 365.94 449.73 ;
   RECT 0.0 449.73 365.94 451.44 ;
   RECT 0.0 451.44 365.94 453.15 ;
   RECT 0.0 453.15 365.94 454.86 ;
   RECT 0.0 454.86 365.94 456.57 ;
   RECT 0.0 456.57 365.94 458.28 ;
   RECT 0.0 458.28 365.94 459.99 ;
   RECT 0.0 459.99 365.94 461.7 ;
   RECT 0.0 461.7 365.94 463.41 ;
   RECT 0.0 463.41 365.94 465.12 ;
   RECT 0.0 465.12 365.94 466.83 ;
   RECT 0.0 466.83 365.94 468.54 ;
   RECT 0.0 468.54 365.94 470.25 ;
   RECT 0.0 470.25 365.94 471.96 ;
   RECT 0.0 471.96 365.94 473.67 ;
   RECT 0.0 473.67 365.94 475.38 ;
  LAYER metal3 ;
   RECT 0.0 0.0 365.94 1.71 ;
   RECT 0.0 1.71 365.94 3.42 ;
   RECT 0.0 3.42 365.94 5.13 ;
   RECT 0.0 5.13 365.94 6.84 ;
   RECT 0.0 6.84 365.94 8.55 ;
   RECT 0.0 8.55 365.94 10.26 ;
   RECT 0.0 10.26 365.94 11.97 ;
   RECT 0.0 11.97 365.94 13.68 ;
   RECT 0.0 13.68 365.94 15.39 ;
   RECT 0.0 15.39 365.94 17.1 ;
   RECT 0.0 17.1 365.94 18.81 ;
   RECT 0.0 18.81 365.94 20.52 ;
   RECT 0.0 20.52 365.94 22.23 ;
   RECT 0.0 22.23 365.94 23.94 ;
   RECT 0.0 23.94 365.94 25.65 ;
   RECT 0.0 25.65 365.94 27.36 ;
   RECT 0.0 27.36 365.94 29.07 ;
   RECT 0.0 29.07 365.94 30.78 ;
   RECT 0.0 30.78 365.94 32.49 ;
   RECT 0.0 32.49 365.94 34.2 ;
   RECT 0.0 34.2 365.94 35.91 ;
   RECT 0.0 35.91 365.94 37.62 ;
   RECT 0.0 37.62 365.94 39.33 ;
   RECT 0.0 39.33 365.94 41.04 ;
   RECT 0.0 41.04 365.94 42.75 ;
   RECT 0.0 42.75 365.94 44.46 ;
   RECT 0.0 44.46 365.94 46.17 ;
   RECT 0.0 46.17 365.94 47.88 ;
   RECT 0.0 47.88 365.94 49.59 ;
   RECT 0.0 49.59 365.94 51.3 ;
   RECT 0.0 51.3 365.94 53.01 ;
   RECT 0.0 53.01 365.94 54.72 ;
   RECT 0.0 54.72 365.94 56.43 ;
   RECT 0.0 56.43 365.94 58.14 ;
   RECT 0.0 58.14 365.94 59.85 ;
   RECT 0.0 59.85 365.94 61.56 ;
   RECT 0.0 61.56 365.94 63.27 ;
   RECT 0.0 63.27 365.94 64.98 ;
   RECT 0.0 64.98 365.94 66.69 ;
   RECT 0.0 66.69 365.94 68.4 ;
   RECT 0.0 68.4 365.94 70.11 ;
   RECT 0.0 70.11 365.94 71.82 ;
   RECT 0.0 71.82 365.94 73.53 ;
   RECT 0.0 73.53 365.94 75.24 ;
   RECT 0.0 75.24 365.94 76.95 ;
   RECT 0.0 76.95 365.94 78.66 ;
   RECT 0.0 78.66 365.94 80.37 ;
   RECT 0.0 80.37 365.94 82.08 ;
   RECT 0.0 82.08 365.94 83.79 ;
   RECT 0.0 83.79 365.94 85.5 ;
   RECT 0.0 85.5 365.94 87.21 ;
   RECT 0.0 87.21 365.94 88.92 ;
   RECT 0.0 88.92 365.94 90.63 ;
   RECT 0.0 90.63 365.94 92.34 ;
   RECT 0.0 92.34 365.94 94.05 ;
   RECT 0.0 94.05 365.94 95.76 ;
   RECT 0.0 95.76 365.94 97.47 ;
   RECT 0.0 97.47 365.94 99.18 ;
   RECT 0.0 99.18 365.94 100.89 ;
   RECT 0.0 100.89 365.94 102.6 ;
   RECT 0.0 102.6 365.94 104.31 ;
   RECT 0.0 104.31 365.94 106.02 ;
   RECT 0.0 106.02 365.94 107.73 ;
   RECT 0.0 107.73 365.94 109.44 ;
   RECT 0.0 109.44 365.94 111.15 ;
   RECT 0.0 111.15 365.94 112.86 ;
   RECT 0.0 112.86 365.94 114.57 ;
   RECT 0.0 114.57 365.94 116.28 ;
   RECT 0.0 116.28 365.94 117.99 ;
   RECT 0.0 117.99 365.94 119.7 ;
   RECT 0.0 119.7 365.94 121.41 ;
   RECT 0.0 121.41 365.94 123.12 ;
   RECT 0.0 123.12 365.94 124.83 ;
   RECT 0.0 124.83 365.94 126.54 ;
   RECT 0.0 126.54 365.94 128.25 ;
   RECT 0.0 128.25 365.94 129.96 ;
   RECT 0.0 129.96 365.94 131.67 ;
   RECT 0.0 131.67 365.94 133.38 ;
   RECT 0.0 133.38 365.94 135.09 ;
   RECT 0.0 135.09 365.94 136.8 ;
   RECT 0.0 136.8 365.94 138.51 ;
   RECT 0.0 138.51 365.94 140.22 ;
   RECT 0.0 140.22 365.94 141.93 ;
   RECT 0.0 141.93 365.94 143.64 ;
   RECT 0.0 143.64 365.94 145.35 ;
   RECT 0.0 145.35 365.94 147.06 ;
   RECT 0.0 147.06 365.94 148.77 ;
   RECT 0.0 148.77 365.94 150.48 ;
   RECT 0.0 150.48 365.94 152.19 ;
   RECT 0.0 152.19 365.94 153.9 ;
   RECT 0.0 153.9 365.94 155.61 ;
   RECT 0.0 155.61 365.94 157.32 ;
   RECT 0.0 157.32 365.94 159.03 ;
   RECT 0.0 159.03 365.94 160.74 ;
   RECT 0.0 160.74 365.94 162.45 ;
   RECT 0.0 162.45 365.94 164.16 ;
   RECT 0.0 164.16 365.94 165.87 ;
   RECT 0.0 165.87 365.94 167.58 ;
   RECT 0.0 167.58 365.94 169.29 ;
   RECT 0.0 169.29 365.94 171.0 ;
   RECT 0.0 171.0 365.94 172.71 ;
   RECT 0.0 172.71 365.94 174.42 ;
   RECT 0.0 174.42 365.94 176.13 ;
   RECT 0.0 176.13 365.94 177.84 ;
   RECT 0.0 177.84 365.94 179.55 ;
   RECT 0.0 179.55 365.94 181.26 ;
   RECT 0.0 181.26 365.94 182.97 ;
   RECT 0.0 182.97 365.94 184.68 ;
   RECT 0.0 184.68 365.94 186.39 ;
   RECT 0.0 186.39 365.94 188.1 ;
   RECT 0.0 188.1 365.94 189.81 ;
   RECT 0.0 189.81 365.94 191.52 ;
   RECT 0.0 191.52 365.94 193.23 ;
   RECT 0.0 193.23 365.94 194.94 ;
   RECT 0.0 194.94 365.94 196.65 ;
   RECT 0.0 196.65 365.94 198.36 ;
   RECT 0.0 198.36 365.94 200.07 ;
   RECT 0.0 200.07 365.94 201.78 ;
   RECT 0.0 201.78 365.94 203.49 ;
   RECT 0.0 203.49 365.94 205.2 ;
   RECT 0.0 205.2 365.94 206.91 ;
   RECT 0.0 206.91 365.94 208.62 ;
   RECT 0.0 208.62 365.94 210.33 ;
   RECT 0.0 210.33 365.94 212.04 ;
   RECT 0.0 212.04 365.94 213.75 ;
   RECT 0.0 213.75 365.94 215.46 ;
   RECT 0.0 215.46 365.94 217.17 ;
   RECT 0.0 217.17 365.94 218.88 ;
   RECT 0.0 218.88 365.94 220.59 ;
   RECT 0.0 220.59 365.94 222.3 ;
   RECT 0.0 222.3 365.94 224.01 ;
   RECT 0.0 224.01 365.94 225.72 ;
   RECT 0.0 225.72 365.94 227.43 ;
   RECT 0.0 227.43 365.94 229.14 ;
   RECT 0.0 229.14 365.94 230.85 ;
   RECT 0.0 230.85 389.12 232.56 ;
   RECT 0.0 232.56 389.12 234.27 ;
   RECT 0.0 234.27 389.12 235.98 ;
   RECT 0.0 235.98 389.12 237.69 ;
   RECT 0.0 237.69 389.12 239.4 ;
   RECT 0.0 239.4 389.12 241.11 ;
   RECT 0.0 241.11 389.12 242.82 ;
   RECT 0.0 242.82 389.12 244.53 ;
   RECT 0.0 244.53 389.12 246.24 ;
   RECT 0.0 246.24 389.12 247.95 ;
   RECT 0.0 247.95 389.12 249.66 ;
   RECT 0.0 249.66 389.12 251.37 ;
   RECT 0.0 251.37 389.12 253.08 ;
   RECT 0.0 253.08 389.12 254.79 ;
   RECT 0.0 254.79 389.12 256.5 ;
   RECT 0.0 256.5 389.12 258.21 ;
   RECT 0.0 258.21 389.12 259.92 ;
   RECT 0.0 259.92 365.94 261.63 ;
   RECT 0.0 261.63 365.94 263.34 ;
   RECT 0.0 263.34 365.94 265.05 ;
   RECT 0.0 265.05 365.94 266.76 ;
   RECT 0.0 266.76 365.94 268.47 ;
   RECT 0.0 268.47 365.94 270.18 ;
   RECT 0.0 270.18 365.94 271.89 ;
   RECT 0.0 271.89 365.94 273.6 ;
   RECT 0.0 273.6 365.94 275.31 ;
   RECT 0.0 275.31 365.94 277.02 ;
   RECT 0.0 277.02 365.94 278.73 ;
   RECT 0.0 278.73 365.94 280.44 ;
   RECT 0.0 280.44 365.94 282.15 ;
   RECT 0.0 282.15 365.94 283.86 ;
   RECT 0.0 283.86 365.94 285.57 ;
   RECT 0.0 285.57 365.94 287.28 ;
   RECT 0.0 287.28 365.94 288.99 ;
   RECT 0.0 288.99 365.94 290.7 ;
   RECT 0.0 290.7 365.94 292.41 ;
   RECT 0.0 292.41 365.94 294.12 ;
   RECT 0.0 294.12 365.94 295.83 ;
   RECT 0.0 295.83 365.94 297.54 ;
   RECT 0.0 297.54 365.94 299.25 ;
   RECT 0.0 299.25 365.94 300.96 ;
   RECT 0.0 300.96 365.94 302.67 ;
   RECT 0.0 302.67 365.94 304.38 ;
   RECT 0.0 304.38 365.94 306.09 ;
   RECT 0.0 306.09 365.94 307.8 ;
   RECT 0.0 307.8 365.94 309.51 ;
   RECT 0.0 309.51 365.94 311.22 ;
   RECT 0.0 311.22 365.94 312.93 ;
   RECT 0.0 312.93 365.94 314.64 ;
   RECT 0.0 314.64 365.94 316.35 ;
   RECT 0.0 316.35 365.94 318.06 ;
   RECT 0.0 318.06 365.94 319.77 ;
   RECT 0.0 319.77 365.94 321.48 ;
   RECT 0.0 321.48 365.94 323.19 ;
   RECT 0.0 323.19 365.94 324.9 ;
   RECT 0.0 324.9 365.94 326.61 ;
   RECT 0.0 326.61 365.94 328.32 ;
   RECT 0.0 328.32 365.94 330.03 ;
   RECT 0.0 330.03 365.94 331.74 ;
   RECT 0.0 331.74 365.94 333.45 ;
   RECT 0.0 333.45 365.94 335.16 ;
   RECT 0.0 335.16 365.94 336.87 ;
   RECT 0.0 336.87 365.94 338.58 ;
   RECT 0.0 338.58 365.94 340.29 ;
   RECT 0.0 340.29 365.94 342.0 ;
   RECT 0.0 342.0 365.94 343.71 ;
   RECT 0.0 343.71 365.94 345.42 ;
   RECT 0.0 345.42 365.94 347.13 ;
   RECT 0.0 347.13 365.94 348.84 ;
   RECT 0.0 348.84 365.94 350.55 ;
   RECT 0.0 350.55 365.94 352.26 ;
   RECT 0.0 352.26 365.94 353.97 ;
   RECT 0.0 353.97 365.94 355.68 ;
   RECT 0.0 355.68 365.94 357.39 ;
   RECT 0.0 357.39 365.94 359.1 ;
   RECT 0.0 359.1 365.94 360.81 ;
   RECT 0.0 360.81 365.94 362.52 ;
   RECT 0.0 362.52 365.94 364.23 ;
   RECT 0.0 364.23 365.94 365.94 ;
   RECT 0.0 365.94 365.94 367.65 ;
   RECT 0.0 367.65 365.94 369.36 ;
   RECT 0.0 369.36 365.94 371.07 ;
   RECT 0.0 371.07 365.94 372.78 ;
   RECT 0.0 372.78 365.94 374.49 ;
   RECT 0.0 374.49 365.94 376.2 ;
   RECT 0.0 376.2 365.94 377.91 ;
   RECT 0.0 377.91 365.94 379.62 ;
   RECT 0.0 379.62 365.94 381.33 ;
   RECT 0.0 381.33 365.94 383.04 ;
   RECT 0.0 383.04 365.94 384.75 ;
   RECT 0.0 384.75 365.94 386.46 ;
   RECT 0.0 386.46 365.94 388.17 ;
   RECT 0.0 388.17 365.94 389.88 ;
   RECT 0.0 389.88 365.94 391.59 ;
   RECT 0.0 391.59 365.94 393.3 ;
   RECT 0.0 393.3 365.94 395.01 ;
   RECT 0.0 395.01 365.94 396.72 ;
   RECT 0.0 396.72 365.94 398.43 ;
   RECT 0.0 398.43 365.94 400.14 ;
   RECT 0.0 400.14 365.94 401.85 ;
   RECT 0.0 401.85 365.94 403.56 ;
   RECT 0.0 403.56 365.94 405.27 ;
   RECT 0.0 405.27 365.94 406.98 ;
   RECT 0.0 406.98 365.94 408.69 ;
   RECT 0.0 408.69 365.94 410.4 ;
   RECT 0.0 410.4 365.94 412.11 ;
   RECT 0.0 412.11 365.94 413.82 ;
   RECT 0.0 413.82 365.94 415.53 ;
   RECT 0.0 415.53 365.94 417.24 ;
   RECT 0.0 417.24 365.94 418.95 ;
   RECT 0.0 418.95 365.94 420.66 ;
   RECT 0.0 420.66 365.94 422.37 ;
   RECT 0.0 422.37 365.94 424.08 ;
   RECT 0.0 424.08 365.94 425.79 ;
   RECT 0.0 425.79 365.94 427.5 ;
   RECT 0.0 427.5 365.94 429.21 ;
   RECT 0.0 429.21 365.94 430.92 ;
   RECT 0.0 430.92 365.94 432.63 ;
   RECT 0.0 432.63 365.94 434.34 ;
   RECT 0.0 434.34 365.94 436.05 ;
   RECT 0.0 436.05 365.94 437.76 ;
   RECT 0.0 437.76 365.94 439.47 ;
   RECT 0.0 439.47 365.94 441.18 ;
   RECT 0.0 441.18 365.94 442.89 ;
   RECT 0.0 442.89 365.94 444.6 ;
   RECT 0.0 444.6 365.94 446.31 ;
   RECT 0.0 446.31 365.94 448.02 ;
   RECT 0.0 448.02 365.94 449.73 ;
   RECT 0.0 449.73 365.94 451.44 ;
   RECT 0.0 451.44 365.94 453.15 ;
   RECT 0.0 453.15 365.94 454.86 ;
   RECT 0.0 454.86 365.94 456.57 ;
   RECT 0.0 456.57 365.94 458.28 ;
   RECT 0.0 458.28 365.94 459.99 ;
   RECT 0.0 459.99 365.94 461.7 ;
   RECT 0.0 461.7 365.94 463.41 ;
   RECT 0.0 463.41 365.94 465.12 ;
   RECT 0.0 465.12 365.94 466.83 ;
   RECT 0.0 466.83 365.94 468.54 ;
   RECT 0.0 468.54 365.94 470.25 ;
   RECT 0.0 470.25 365.94 471.96 ;
   RECT 0.0 471.96 365.94 473.67 ;
   RECT 0.0 473.67 365.94 475.38 ;
  LAYER via3 ;
   RECT 0.0 0.0 365.94 1.71 ;
   RECT 0.0 1.71 365.94 3.42 ;
   RECT 0.0 3.42 365.94 5.13 ;
   RECT 0.0 5.13 365.94 6.84 ;
   RECT 0.0 6.84 365.94 8.55 ;
   RECT 0.0 8.55 365.94 10.26 ;
   RECT 0.0 10.26 365.94 11.97 ;
   RECT 0.0 11.97 365.94 13.68 ;
   RECT 0.0 13.68 365.94 15.39 ;
   RECT 0.0 15.39 365.94 17.1 ;
   RECT 0.0 17.1 365.94 18.81 ;
   RECT 0.0 18.81 365.94 20.52 ;
   RECT 0.0 20.52 365.94 22.23 ;
   RECT 0.0 22.23 365.94 23.94 ;
   RECT 0.0 23.94 365.94 25.65 ;
   RECT 0.0 25.65 365.94 27.36 ;
   RECT 0.0 27.36 365.94 29.07 ;
   RECT 0.0 29.07 365.94 30.78 ;
   RECT 0.0 30.78 365.94 32.49 ;
   RECT 0.0 32.49 365.94 34.2 ;
   RECT 0.0 34.2 365.94 35.91 ;
   RECT 0.0 35.91 365.94 37.62 ;
   RECT 0.0 37.62 365.94 39.33 ;
   RECT 0.0 39.33 365.94 41.04 ;
   RECT 0.0 41.04 365.94 42.75 ;
   RECT 0.0 42.75 365.94 44.46 ;
   RECT 0.0 44.46 365.94 46.17 ;
   RECT 0.0 46.17 365.94 47.88 ;
   RECT 0.0 47.88 365.94 49.59 ;
   RECT 0.0 49.59 365.94 51.3 ;
   RECT 0.0 51.3 365.94 53.01 ;
   RECT 0.0 53.01 365.94 54.72 ;
   RECT 0.0 54.72 365.94 56.43 ;
   RECT 0.0 56.43 365.94 58.14 ;
   RECT 0.0 58.14 365.94 59.85 ;
   RECT 0.0 59.85 365.94 61.56 ;
   RECT 0.0 61.56 365.94 63.27 ;
   RECT 0.0 63.27 365.94 64.98 ;
   RECT 0.0 64.98 365.94 66.69 ;
   RECT 0.0 66.69 365.94 68.4 ;
   RECT 0.0 68.4 365.94 70.11 ;
   RECT 0.0 70.11 365.94 71.82 ;
   RECT 0.0 71.82 365.94 73.53 ;
   RECT 0.0 73.53 365.94 75.24 ;
   RECT 0.0 75.24 365.94 76.95 ;
   RECT 0.0 76.95 365.94 78.66 ;
   RECT 0.0 78.66 365.94 80.37 ;
   RECT 0.0 80.37 365.94 82.08 ;
   RECT 0.0 82.08 365.94 83.79 ;
   RECT 0.0 83.79 365.94 85.5 ;
   RECT 0.0 85.5 365.94 87.21 ;
   RECT 0.0 87.21 365.94 88.92 ;
   RECT 0.0 88.92 365.94 90.63 ;
   RECT 0.0 90.63 365.94 92.34 ;
   RECT 0.0 92.34 365.94 94.05 ;
   RECT 0.0 94.05 365.94 95.76 ;
   RECT 0.0 95.76 365.94 97.47 ;
   RECT 0.0 97.47 365.94 99.18 ;
   RECT 0.0 99.18 365.94 100.89 ;
   RECT 0.0 100.89 365.94 102.6 ;
   RECT 0.0 102.6 365.94 104.31 ;
   RECT 0.0 104.31 365.94 106.02 ;
   RECT 0.0 106.02 365.94 107.73 ;
   RECT 0.0 107.73 365.94 109.44 ;
   RECT 0.0 109.44 365.94 111.15 ;
   RECT 0.0 111.15 365.94 112.86 ;
   RECT 0.0 112.86 365.94 114.57 ;
   RECT 0.0 114.57 365.94 116.28 ;
   RECT 0.0 116.28 365.94 117.99 ;
   RECT 0.0 117.99 365.94 119.7 ;
   RECT 0.0 119.7 365.94 121.41 ;
   RECT 0.0 121.41 365.94 123.12 ;
   RECT 0.0 123.12 365.94 124.83 ;
   RECT 0.0 124.83 365.94 126.54 ;
   RECT 0.0 126.54 365.94 128.25 ;
   RECT 0.0 128.25 365.94 129.96 ;
   RECT 0.0 129.96 365.94 131.67 ;
   RECT 0.0 131.67 365.94 133.38 ;
   RECT 0.0 133.38 365.94 135.09 ;
   RECT 0.0 135.09 365.94 136.8 ;
   RECT 0.0 136.8 365.94 138.51 ;
   RECT 0.0 138.51 365.94 140.22 ;
   RECT 0.0 140.22 365.94 141.93 ;
   RECT 0.0 141.93 365.94 143.64 ;
   RECT 0.0 143.64 365.94 145.35 ;
   RECT 0.0 145.35 365.94 147.06 ;
   RECT 0.0 147.06 365.94 148.77 ;
   RECT 0.0 148.77 365.94 150.48 ;
   RECT 0.0 150.48 365.94 152.19 ;
   RECT 0.0 152.19 365.94 153.9 ;
   RECT 0.0 153.9 365.94 155.61 ;
   RECT 0.0 155.61 365.94 157.32 ;
   RECT 0.0 157.32 365.94 159.03 ;
   RECT 0.0 159.03 365.94 160.74 ;
   RECT 0.0 160.74 365.94 162.45 ;
   RECT 0.0 162.45 365.94 164.16 ;
   RECT 0.0 164.16 365.94 165.87 ;
   RECT 0.0 165.87 365.94 167.58 ;
   RECT 0.0 167.58 365.94 169.29 ;
   RECT 0.0 169.29 365.94 171.0 ;
   RECT 0.0 171.0 365.94 172.71 ;
   RECT 0.0 172.71 365.94 174.42 ;
   RECT 0.0 174.42 365.94 176.13 ;
   RECT 0.0 176.13 365.94 177.84 ;
   RECT 0.0 177.84 365.94 179.55 ;
   RECT 0.0 179.55 365.94 181.26 ;
   RECT 0.0 181.26 365.94 182.97 ;
   RECT 0.0 182.97 365.94 184.68 ;
   RECT 0.0 184.68 365.94 186.39 ;
   RECT 0.0 186.39 365.94 188.1 ;
   RECT 0.0 188.1 365.94 189.81 ;
   RECT 0.0 189.81 365.94 191.52 ;
   RECT 0.0 191.52 365.94 193.23 ;
   RECT 0.0 193.23 365.94 194.94 ;
   RECT 0.0 194.94 365.94 196.65 ;
   RECT 0.0 196.65 365.94 198.36 ;
   RECT 0.0 198.36 365.94 200.07 ;
   RECT 0.0 200.07 365.94 201.78 ;
   RECT 0.0 201.78 365.94 203.49 ;
   RECT 0.0 203.49 365.94 205.2 ;
   RECT 0.0 205.2 365.94 206.91 ;
   RECT 0.0 206.91 365.94 208.62 ;
   RECT 0.0 208.62 365.94 210.33 ;
   RECT 0.0 210.33 365.94 212.04 ;
   RECT 0.0 212.04 365.94 213.75 ;
   RECT 0.0 213.75 365.94 215.46 ;
   RECT 0.0 215.46 365.94 217.17 ;
   RECT 0.0 217.17 365.94 218.88 ;
   RECT 0.0 218.88 365.94 220.59 ;
   RECT 0.0 220.59 365.94 222.3 ;
   RECT 0.0 222.3 365.94 224.01 ;
   RECT 0.0 224.01 365.94 225.72 ;
   RECT 0.0 225.72 365.94 227.43 ;
   RECT 0.0 227.43 365.94 229.14 ;
   RECT 0.0 229.14 365.94 230.85 ;
   RECT 0.0 230.85 389.12 232.56 ;
   RECT 0.0 232.56 389.12 234.27 ;
   RECT 0.0 234.27 389.12 235.98 ;
   RECT 0.0 235.98 389.12 237.69 ;
   RECT 0.0 237.69 389.12 239.4 ;
   RECT 0.0 239.4 389.12 241.11 ;
   RECT 0.0 241.11 389.12 242.82 ;
   RECT 0.0 242.82 389.12 244.53 ;
   RECT 0.0 244.53 389.12 246.24 ;
   RECT 0.0 246.24 389.12 247.95 ;
   RECT 0.0 247.95 389.12 249.66 ;
   RECT 0.0 249.66 389.12 251.37 ;
   RECT 0.0 251.37 389.12 253.08 ;
   RECT 0.0 253.08 389.12 254.79 ;
   RECT 0.0 254.79 389.12 256.5 ;
   RECT 0.0 256.5 389.12 258.21 ;
   RECT 0.0 258.21 389.12 259.92 ;
   RECT 0.0 259.92 365.94 261.63 ;
   RECT 0.0 261.63 365.94 263.34 ;
   RECT 0.0 263.34 365.94 265.05 ;
   RECT 0.0 265.05 365.94 266.76 ;
   RECT 0.0 266.76 365.94 268.47 ;
   RECT 0.0 268.47 365.94 270.18 ;
   RECT 0.0 270.18 365.94 271.89 ;
   RECT 0.0 271.89 365.94 273.6 ;
   RECT 0.0 273.6 365.94 275.31 ;
   RECT 0.0 275.31 365.94 277.02 ;
   RECT 0.0 277.02 365.94 278.73 ;
   RECT 0.0 278.73 365.94 280.44 ;
   RECT 0.0 280.44 365.94 282.15 ;
   RECT 0.0 282.15 365.94 283.86 ;
   RECT 0.0 283.86 365.94 285.57 ;
   RECT 0.0 285.57 365.94 287.28 ;
   RECT 0.0 287.28 365.94 288.99 ;
   RECT 0.0 288.99 365.94 290.7 ;
   RECT 0.0 290.7 365.94 292.41 ;
   RECT 0.0 292.41 365.94 294.12 ;
   RECT 0.0 294.12 365.94 295.83 ;
   RECT 0.0 295.83 365.94 297.54 ;
   RECT 0.0 297.54 365.94 299.25 ;
   RECT 0.0 299.25 365.94 300.96 ;
   RECT 0.0 300.96 365.94 302.67 ;
   RECT 0.0 302.67 365.94 304.38 ;
   RECT 0.0 304.38 365.94 306.09 ;
   RECT 0.0 306.09 365.94 307.8 ;
   RECT 0.0 307.8 365.94 309.51 ;
   RECT 0.0 309.51 365.94 311.22 ;
   RECT 0.0 311.22 365.94 312.93 ;
   RECT 0.0 312.93 365.94 314.64 ;
   RECT 0.0 314.64 365.94 316.35 ;
   RECT 0.0 316.35 365.94 318.06 ;
   RECT 0.0 318.06 365.94 319.77 ;
   RECT 0.0 319.77 365.94 321.48 ;
   RECT 0.0 321.48 365.94 323.19 ;
   RECT 0.0 323.19 365.94 324.9 ;
   RECT 0.0 324.9 365.94 326.61 ;
   RECT 0.0 326.61 365.94 328.32 ;
   RECT 0.0 328.32 365.94 330.03 ;
   RECT 0.0 330.03 365.94 331.74 ;
   RECT 0.0 331.74 365.94 333.45 ;
   RECT 0.0 333.45 365.94 335.16 ;
   RECT 0.0 335.16 365.94 336.87 ;
   RECT 0.0 336.87 365.94 338.58 ;
   RECT 0.0 338.58 365.94 340.29 ;
   RECT 0.0 340.29 365.94 342.0 ;
   RECT 0.0 342.0 365.94 343.71 ;
   RECT 0.0 343.71 365.94 345.42 ;
   RECT 0.0 345.42 365.94 347.13 ;
   RECT 0.0 347.13 365.94 348.84 ;
   RECT 0.0 348.84 365.94 350.55 ;
   RECT 0.0 350.55 365.94 352.26 ;
   RECT 0.0 352.26 365.94 353.97 ;
   RECT 0.0 353.97 365.94 355.68 ;
   RECT 0.0 355.68 365.94 357.39 ;
   RECT 0.0 357.39 365.94 359.1 ;
   RECT 0.0 359.1 365.94 360.81 ;
   RECT 0.0 360.81 365.94 362.52 ;
   RECT 0.0 362.52 365.94 364.23 ;
   RECT 0.0 364.23 365.94 365.94 ;
   RECT 0.0 365.94 365.94 367.65 ;
   RECT 0.0 367.65 365.94 369.36 ;
   RECT 0.0 369.36 365.94 371.07 ;
   RECT 0.0 371.07 365.94 372.78 ;
   RECT 0.0 372.78 365.94 374.49 ;
   RECT 0.0 374.49 365.94 376.2 ;
   RECT 0.0 376.2 365.94 377.91 ;
   RECT 0.0 377.91 365.94 379.62 ;
   RECT 0.0 379.62 365.94 381.33 ;
   RECT 0.0 381.33 365.94 383.04 ;
   RECT 0.0 383.04 365.94 384.75 ;
   RECT 0.0 384.75 365.94 386.46 ;
   RECT 0.0 386.46 365.94 388.17 ;
   RECT 0.0 388.17 365.94 389.88 ;
   RECT 0.0 389.88 365.94 391.59 ;
   RECT 0.0 391.59 365.94 393.3 ;
   RECT 0.0 393.3 365.94 395.01 ;
   RECT 0.0 395.01 365.94 396.72 ;
   RECT 0.0 396.72 365.94 398.43 ;
   RECT 0.0 398.43 365.94 400.14 ;
   RECT 0.0 400.14 365.94 401.85 ;
   RECT 0.0 401.85 365.94 403.56 ;
   RECT 0.0 403.56 365.94 405.27 ;
   RECT 0.0 405.27 365.94 406.98 ;
   RECT 0.0 406.98 365.94 408.69 ;
   RECT 0.0 408.69 365.94 410.4 ;
   RECT 0.0 410.4 365.94 412.11 ;
   RECT 0.0 412.11 365.94 413.82 ;
   RECT 0.0 413.82 365.94 415.53 ;
   RECT 0.0 415.53 365.94 417.24 ;
   RECT 0.0 417.24 365.94 418.95 ;
   RECT 0.0 418.95 365.94 420.66 ;
   RECT 0.0 420.66 365.94 422.37 ;
   RECT 0.0 422.37 365.94 424.08 ;
   RECT 0.0 424.08 365.94 425.79 ;
   RECT 0.0 425.79 365.94 427.5 ;
   RECT 0.0 427.5 365.94 429.21 ;
   RECT 0.0 429.21 365.94 430.92 ;
   RECT 0.0 430.92 365.94 432.63 ;
   RECT 0.0 432.63 365.94 434.34 ;
   RECT 0.0 434.34 365.94 436.05 ;
   RECT 0.0 436.05 365.94 437.76 ;
   RECT 0.0 437.76 365.94 439.47 ;
   RECT 0.0 439.47 365.94 441.18 ;
   RECT 0.0 441.18 365.94 442.89 ;
   RECT 0.0 442.89 365.94 444.6 ;
   RECT 0.0 444.6 365.94 446.31 ;
   RECT 0.0 446.31 365.94 448.02 ;
   RECT 0.0 448.02 365.94 449.73 ;
   RECT 0.0 449.73 365.94 451.44 ;
   RECT 0.0 451.44 365.94 453.15 ;
   RECT 0.0 453.15 365.94 454.86 ;
   RECT 0.0 454.86 365.94 456.57 ;
   RECT 0.0 456.57 365.94 458.28 ;
   RECT 0.0 458.28 365.94 459.99 ;
   RECT 0.0 459.99 365.94 461.7 ;
   RECT 0.0 461.7 365.94 463.41 ;
   RECT 0.0 463.41 365.94 465.12 ;
   RECT 0.0 465.12 365.94 466.83 ;
   RECT 0.0 466.83 365.94 468.54 ;
   RECT 0.0 468.54 365.94 470.25 ;
   RECT 0.0 470.25 365.94 471.96 ;
   RECT 0.0 471.96 365.94 473.67 ;
   RECT 0.0 473.67 365.94 475.38 ;
  LAYER metal4 ;
   RECT 0.0 0.0 365.94 1.71 ;
   RECT 0.0 1.71 365.94 3.42 ;
   RECT 0.0 3.42 365.94 5.13 ;
   RECT 0.0 5.13 365.94 6.84 ;
   RECT 0.0 6.84 365.94 8.55 ;
   RECT 0.0 8.55 365.94 10.26 ;
   RECT 0.0 10.26 365.94 11.97 ;
   RECT 0.0 11.97 365.94 13.68 ;
   RECT 0.0 13.68 365.94 15.39 ;
   RECT 0.0 15.39 365.94 17.1 ;
   RECT 0.0 17.1 365.94 18.81 ;
   RECT 0.0 18.81 365.94 20.52 ;
   RECT 0.0 20.52 365.94 22.23 ;
   RECT 0.0 22.23 365.94 23.94 ;
   RECT 0.0 23.94 365.94 25.65 ;
   RECT 0.0 25.65 365.94 27.36 ;
   RECT 0.0 27.36 365.94 29.07 ;
   RECT 0.0 29.07 365.94 30.78 ;
   RECT 0.0 30.78 365.94 32.49 ;
   RECT 0.0 32.49 365.94 34.2 ;
   RECT 0.0 34.2 365.94 35.91 ;
   RECT 0.0 35.91 365.94 37.62 ;
   RECT 0.0 37.62 365.94 39.33 ;
   RECT 0.0 39.33 365.94 41.04 ;
   RECT 0.0 41.04 365.94 42.75 ;
   RECT 0.0 42.75 365.94 44.46 ;
   RECT 0.0 44.46 365.94 46.17 ;
   RECT 0.0 46.17 365.94 47.88 ;
   RECT 0.0 47.88 365.94 49.59 ;
   RECT 0.0 49.59 365.94 51.3 ;
   RECT 0.0 51.3 365.94 53.01 ;
   RECT 0.0 53.01 365.94 54.72 ;
   RECT 0.0 54.72 365.94 56.43 ;
   RECT 0.0 56.43 365.94 58.14 ;
   RECT 0.0 58.14 365.94 59.85 ;
   RECT 0.0 59.85 365.94 61.56 ;
   RECT 0.0 61.56 365.94 63.27 ;
   RECT 0.0 63.27 365.94 64.98 ;
   RECT 0.0 64.98 365.94 66.69 ;
   RECT 0.0 66.69 365.94 68.4 ;
   RECT 0.0 68.4 365.94 70.11 ;
   RECT 0.0 70.11 365.94 71.82 ;
   RECT 0.0 71.82 365.94 73.53 ;
   RECT 0.0 73.53 365.94 75.24 ;
   RECT 0.0 75.24 365.94 76.95 ;
   RECT 0.0 76.95 365.94 78.66 ;
   RECT 0.0 78.66 365.94 80.37 ;
   RECT 0.0 80.37 365.94 82.08 ;
   RECT 0.0 82.08 365.94 83.79 ;
   RECT 0.0 83.79 365.94 85.5 ;
   RECT 0.0 85.5 365.94 87.21 ;
   RECT 0.0 87.21 365.94 88.92 ;
   RECT 0.0 88.92 365.94 90.63 ;
   RECT 0.0 90.63 365.94 92.34 ;
   RECT 0.0 92.34 365.94 94.05 ;
   RECT 0.0 94.05 365.94 95.76 ;
   RECT 0.0 95.76 365.94 97.47 ;
   RECT 0.0 97.47 365.94 99.18 ;
   RECT 0.0 99.18 365.94 100.89 ;
   RECT 0.0 100.89 365.94 102.6 ;
   RECT 0.0 102.6 365.94 104.31 ;
   RECT 0.0 104.31 365.94 106.02 ;
   RECT 0.0 106.02 365.94 107.73 ;
   RECT 0.0 107.73 365.94 109.44 ;
   RECT 0.0 109.44 365.94 111.15 ;
   RECT 0.0 111.15 365.94 112.86 ;
   RECT 0.0 112.86 365.94 114.57 ;
   RECT 0.0 114.57 365.94 116.28 ;
   RECT 0.0 116.28 365.94 117.99 ;
   RECT 0.0 117.99 365.94 119.7 ;
   RECT 0.0 119.7 365.94 121.41 ;
   RECT 0.0 121.41 365.94 123.12 ;
   RECT 0.0 123.12 365.94 124.83 ;
   RECT 0.0 124.83 365.94 126.54 ;
   RECT 0.0 126.54 365.94 128.25 ;
   RECT 0.0 128.25 365.94 129.96 ;
   RECT 0.0 129.96 365.94 131.67 ;
   RECT 0.0 131.67 365.94 133.38 ;
   RECT 0.0 133.38 365.94 135.09 ;
   RECT 0.0 135.09 365.94 136.8 ;
   RECT 0.0 136.8 365.94 138.51 ;
   RECT 0.0 138.51 365.94 140.22 ;
   RECT 0.0 140.22 365.94 141.93 ;
   RECT 0.0 141.93 365.94 143.64 ;
   RECT 0.0 143.64 365.94 145.35 ;
   RECT 0.0 145.35 365.94 147.06 ;
   RECT 0.0 147.06 365.94 148.77 ;
   RECT 0.0 148.77 365.94 150.48 ;
   RECT 0.0 150.48 365.94 152.19 ;
   RECT 0.0 152.19 365.94 153.9 ;
   RECT 0.0 153.9 365.94 155.61 ;
   RECT 0.0 155.61 365.94 157.32 ;
   RECT 0.0 157.32 365.94 159.03 ;
   RECT 0.0 159.03 365.94 160.74 ;
   RECT 0.0 160.74 365.94 162.45 ;
   RECT 0.0 162.45 365.94 164.16 ;
   RECT 0.0 164.16 365.94 165.87 ;
   RECT 0.0 165.87 365.94 167.58 ;
   RECT 0.0 167.58 365.94 169.29 ;
   RECT 0.0 169.29 365.94 171.0 ;
   RECT 0.0 171.0 365.94 172.71 ;
   RECT 0.0 172.71 365.94 174.42 ;
   RECT 0.0 174.42 365.94 176.13 ;
   RECT 0.0 176.13 365.94 177.84 ;
   RECT 0.0 177.84 365.94 179.55 ;
   RECT 0.0 179.55 365.94 181.26 ;
   RECT 0.0 181.26 365.94 182.97 ;
   RECT 0.0 182.97 365.94 184.68 ;
   RECT 0.0 184.68 365.94 186.39 ;
   RECT 0.0 186.39 365.94 188.1 ;
   RECT 0.0 188.1 365.94 189.81 ;
   RECT 0.0 189.81 365.94 191.52 ;
   RECT 0.0 191.52 365.94 193.23 ;
   RECT 0.0 193.23 365.94 194.94 ;
   RECT 0.0 194.94 365.94 196.65 ;
   RECT 0.0 196.65 365.94 198.36 ;
   RECT 0.0 198.36 365.94 200.07 ;
   RECT 0.0 200.07 365.94 201.78 ;
   RECT 0.0 201.78 365.94 203.49 ;
   RECT 0.0 203.49 365.94 205.2 ;
   RECT 0.0 205.2 365.94 206.91 ;
   RECT 0.0 206.91 365.94 208.62 ;
   RECT 0.0 208.62 365.94 210.33 ;
   RECT 0.0 210.33 365.94 212.04 ;
   RECT 0.0 212.04 365.94 213.75 ;
   RECT 0.0 213.75 365.94 215.46 ;
   RECT 0.0 215.46 365.94 217.17 ;
   RECT 0.0 217.17 365.94 218.88 ;
   RECT 0.0 218.88 365.94 220.59 ;
   RECT 0.0 220.59 365.94 222.3 ;
   RECT 0.0 222.3 365.94 224.01 ;
   RECT 0.0 224.01 365.94 225.72 ;
   RECT 0.0 225.72 365.94 227.43 ;
   RECT 0.0 227.43 365.94 229.14 ;
   RECT 0.0 229.14 365.94 230.85 ;
   RECT 0.0 230.85 389.12 232.56 ;
   RECT 0.0 232.56 389.12 234.27 ;
   RECT 0.0 234.27 389.12 235.98 ;
   RECT 0.0 235.98 389.12 237.69 ;
   RECT 0.0 237.69 389.12 239.4 ;
   RECT 0.0 239.4 389.12 241.11 ;
   RECT 0.0 241.11 389.12 242.82 ;
   RECT 0.0 242.82 389.12 244.53 ;
   RECT 0.0 244.53 389.12 246.24 ;
   RECT 0.0 246.24 389.12 247.95 ;
   RECT 0.0 247.95 389.12 249.66 ;
   RECT 0.0 249.66 389.12 251.37 ;
   RECT 0.0 251.37 389.12 253.08 ;
   RECT 0.0 253.08 389.12 254.79 ;
   RECT 0.0 254.79 389.12 256.5 ;
   RECT 0.0 256.5 389.12 258.21 ;
   RECT 0.0 258.21 389.12 259.92 ;
   RECT 0.0 259.92 365.94 261.63 ;
   RECT 0.0 261.63 365.94 263.34 ;
   RECT 0.0 263.34 365.94 265.05 ;
   RECT 0.0 265.05 365.94 266.76 ;
   RECT 0.0 266.76 365.94 268.47 ;
   RECT 0.0 268.47 365.94 270.18 ;
   RECT 0.0 270.18 365.94 271.89 ;
   RECT 0.0 271.89 365.94 273.6 ;
   RECT 0.0 273.6 365.94 275.31 ;
   RECT 0.0 275.31 365.94 277.02 ;
   RECT 0.0 277.02 365.94 278.73 ;
   RECT 0.0 278.73 365.94 280.44 ;
   RECT 0.0 280.44 365.94 282.15 ;
   RECT 0.0 282.15 365.94 283.86 ;
   RECT 0.0 283.86 365.94 285.57 ;
   RECT 0.0 285.57 365.94 287.28 ;
   RECT 0.0 287.28 365.94 288.99 ;
   RECT 0.0 288.99 365.94 290.7 ;
   RECT 0.0 290.7 365.94 292.41 ;
   RECT 0.0 292.41 365.94 294.12 ;
   RECT 0.0 294.12 365.94 295.83 ;
   RECT 0.0 295.83 365.94 297.54 ;
   RECT 0.0 297.54 365.94 299.25 ;
   RECT 0.0 299.25 365.94 300.96 ;
   RECT 0.0 300.96 365.94 302.67 ;
   RECT 0.0 302.67 365.94 304.38 ;
   RECT 0.0 304.38 365.94 306.09 ;
   RECT 0.0 306.09 365.94 307.8 ;
   RECT 0.0 307.8 365.94 309.51 ;
   RECT 0.0 309.51 365.94 311.22 ;
   RECT 0.0 311.22 365.94 312.93 ;
   RECT 0.0 312.93 365.94 314.64 ;
   RECT 0.0 314.64 365.94 316.35 ;
   RECT 0.0 316.35 365.94 318.06 ;
   RECT 0.0 318.06 365.94 319.77 ;
   RECT 0.0 319.77 365.94 321.48 ;
   RECT 0.0 321.48 365.94 323.19 ;
   RECT 0.0 323.19 365.94 324.9 ;
   RECT 0.0 324.9 365.94 326.61 ;
   RECT 0.0 326.61 365.94 328.32 ;
   RECT 0.0 328.32 365.94 330.03 ;
   RECT 0.0 330.03 365.94 331.74 ;
   RECT 0.0 331.74 365.94 333.45 ;
   RECT 0.0 333.45 365.94 335.16 ;
   RECT 0.0 335.16 365.94 336.87 ;
   RECT 0.0 336.87 365.94 338.58 ;
   RECT 0.0 338.58 365.94 340.29 ;
   RECT 0.0 340.29 365.94 342.0 ;
   RECT 0.0 342.0 365.94 343.71 ;
   RECT 0.0 343.71 365.94 345.42 ;
   RECT 0.0 345.42 365.94 347.13 ;
   RECT 0.0 347.13 365.94 348.84 ;
   RECT 0.0 348.84 365.94 350.55 ;
   RECT 0.0 350.55 365.94 352.26 ;
   RECT 0.0 352.26 365.94 353.97 ;
   RECT 0.0 353.97 365.94 355.68 ;
   RECT 0.0 355.68 365.94 357.39 ;
   RECT 0.0 357.39 365.94 359.1 ;
   RECT 0.0 359.1 365.94 360.81 ;
   RECT 0.0 360.81 365.94 362.52 ;
   RECT 0.0 362.52 365.94 364.23 ;
   RECT 0.0 364.23 365.94 365.94 ;
   RECT 0.0 365.94 365.94 367.65 ;
   RECT 0.0 367.65 365.94 369.36 ;
   RECT 0.0 369.36 365.94 371.07 ;
   RECT 0.0 371.07 365.94 372.78 ;
   RECT 0.0 372.78 365.94 374.49 ;
   RECT 0.0 374.49 365.94 376.2 ;
   RECT 0.0 376.2 365.94 377.91 ;
   RECT 0.0 377.91 365.94 379.62 ;
   RECT 0.0 379.62 365.94 381.33 ;
   RECT 0.0 381.33 365.94 383.04 ;
   RECT 0.0 383.04 365.94 384.75 ;
   RECT 0.0 384.75 365.94 386.46 ;
   RECT 0.0 386.46 365.94 388.17 ;
   RECT 0.0 388.17 365.94 389.88 ;
   RECT 0.0 389.88 365.94 391.59 ;
   RECT 0.0 391.59 365.94 393.3 ;
   RECT 0.0 393.3 365.94 395.01 ;
   RECT 0.0 395.01 365.94 396.72 ;
   RECT 0.0 396.72 365.94 398.43 ;
   RECT 0.0 398.43 365.94 400.14 ;
   RECT 0.0 400.14 365.94 401.85 ;
   RECT 0.0 401.85 365.94 403.56 ;
   RECT 0.0 403.56 365.94 405.27 ;
   RECT 0.0 405.27 365.94 406.98 ;
   RECT 0.0 406.98 365.94 408.69 ;
   RECT 0.0 408.69 365.94 410.4 ;
   RECT 0.0 410.4 365.94 412.11 ;
   RECT 0.0 412.11 365.94 413.82 ;
   RECT 0.0 413.82 365.94 415.53 ;
   RECT 0.0 415.53 365.94 417.24 ;
   RECT 0.0 417.24 365.94 418.95 ;
   RECT 0.0 418.95 365.94 420.66 ;
   RECT 0.0 420.66 365.94 422.37 ;
   RECT 0.0 422.37 365.94 424.08 ;
   RECT 0.0 424.08 365.94 425.79 ;
   RECT 0.0 425.79 365.94 427.5 ;
   RECT 0.0 427.5 365.94 429.21 ;
   RECT 0.0 429.21 365.94 430.92 ;
   RECT 0.0 430.92 365.94 432.63 ;
   RECT 0.0 432.63 365.94 434.34 ;
   RECT 0.0 434.34 365.94 436.05 ;
   RECT 0.0 436.05 365.94 437.76 ;
   RECT 0.0 437.76 365.94 439.47 ;
   RECT 0.0 439.47 365.94 441.18 ;
   RECT 0.0 441.18 365.94 442.89 ;
   RECT 0.0 442.89 365.94 444.6 ;
   RECT 0.0 444.6 365.94 446.31 ;
   RECT 0.0 446.31 365.94 448.02 ;
   RECT 0.0 448.02 365.94 449.73 ;
   RECT 0.0 449.73 365.94 451.44 ;
   RECT 0.0 451.44 365.94 453.15 ;
   RECT 0.0 453.15 365.94 454.86 ;
   RECT 0.0 454.86 365.94 456.57 ;
   RECT 0.0 456.57 365.94 458.28 ;
   RECT 0.0 458.28 365.94 459.99 ;
   RECT 0.0 459.99 365.94 461.7 ;
   RECT 0.0 461.7 365.94 463.41 ;
   RECT 0.0 463.41 365.94 465.12 ;
   RECT 0.0 465.12 365.94 466.83 ;
   RECT 0.0 466.83 365.94 468.54 ;
   RECT 0.0 468.54 365.94 470.25 ;
   RECT 0.0 470.25 365.94 471.96 ;
   RECT 0.0 471.96 365.94 473.67 ;
   RECT 0.0 473.67 365.94 475.38 ;
 END
END block_1024x2502_161

MACRO block_341x369_82
 CLASS BLOCK ;
 FOREIGN block_341x369_82 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 129.58 BY 70.11 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 20.235 126.445 20.805 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 26.695 126.445 27.265 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 6.935 3.325 7.505 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 6.935 4.085 7.505 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 9.215 3.325 9.785 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 10.735 3.325 11.305 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 11.875 3.325 12.445 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 13.015 3.325 13.585 ;
  END
 END o7
 PIN o8
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 13.395 4.085 13.965 ;
  END
 END o8
 PIN o9
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 13.775 3.325 14.345 ;
  END
 END o9
 PIN o10
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 15.295 3.325 15.865 ;
  END
 END o10
 PIN o11
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 16.055 3.325 16.625 ;
  END
 END o11
 PIN o12
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 16.815 3.325 17.385 ;
  END
 END o12
 PIN o13
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 12.635 4.085 13.205 ;
  END
 END o13
 PIN o14
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 19.855 3.325 20.425 ;
  END
 END o14
 PIN o15
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 20.615 3.325 21.185 ;
  END
 END o15
 PIN o16
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 21.375 3.325 21.945 ;
  END
 END o16
 PIN o17
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 22.135 3.325 22.705 ;
  END
 END o17
 PIN o18
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 22.895 3.325 23.465 ;
  END
 END o18
 PIN o19
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 18.335 3.325 18.905 ;
  END
 END o19
 PIN o20
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 25.935 3.325 26.505 ;
  END
 END o20
 PIN o21
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 26.695 3.325 27.265 ;
  END
 END o21
 PIN o22
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 27.455 3.325 28.025 ;
  END
 END o22
 PIN o23
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 28.975 3.325 29.545 ;
  END
 END o23
 PIN o24
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 29.735 3.325 30.305 ;
  END
 END o24
 PIN o25
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 25.175 3.325 25.745 ;
  END
 END o25
 PIN o26
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 32.015 3.325 32.585 ;
  END
 END o26
 PIN o27
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 33.535 3.325 34.105 ;
  END
 END o27
 PIN o28
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 34.295 3.325 34.865 ;
  END
 END o28
 PIN o29
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 35.055 3.325 35.625 ;
  END
 END o29
 PIN o30
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 35.815 3.325 36.385 ;
  END
 END o30
 PIN o31
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 31.255 3.325 31.825 ;
  END
 END o31
 PIN o32
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 38.095 126.445 38.665 ;
  END
 END o32
 PIN o33
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 38.855 126.445 39.425 ;
  END
 END o33
 PIN o34
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 39.615 126.445 40.185 ;
  END
 END o34
 PIN o35
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 42.655 126.445 43.225 ;
  END
 END o35
 PIN o36
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 29.735 126.445 30.305 ;
  END
 END o36
 PIN o37
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 21.755 126.445 22.325 ;
  END
 END o37
 PIN o38
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 31.255 126.445 31.825 ;
  END
 END o38
 PIN o39
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 32.015 126.445 32.585 ;
  END
 END o39
 PIN o40
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 33.535 126.445 34.105 ;
  END
 END o40
 PIN o41
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 34.295 126.445 34.865 ;
  END
 END o41
 PIN o42
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 35.055 126.445 35.625 ;
  END
 END o42
 PIN o43
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 30.495 126.445 31.065 ;
  END
 END o43
 PIN o44
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 28.975 126.445 29.545 ;
  END
 END o44
 PIN o45
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 41.135 3.325 41.705 ;
  END
 END o45
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 35.815 126.445 36.385 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 43.035 125.685 43.605 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 32.395 125.685 32.965 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 35.435 125.685 36.005 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 36.955 126.445 37.525 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 36.575 125.685 37.145 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 33.915 125.685 34.485 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 30.115 125.685 30.685 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 40.375 3.325 40.945 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 8.455 3.325 9.025 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 25.935 126.445 26.505 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 25.175 126.445 25.745 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 24.415 126.445 24.985 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 34.675 125.685 35.245 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 30.875 125.685 31.445 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 40.755 126.445 41.325 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 27.455 126.445 28.025 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 38.475 125.685 39.045 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 39.995 125.685 40.565 ;
  END
 END i18
 PIN i19
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 39.235 125.685 39.805 ;
  END
 END i19
 PIN i20
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 124.355 40.375 124.925 40.945 ;
  END
 END i20
 PIN i21
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 8.455 126.445 9.025 ;
  END
 END i21
 PIN i22
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 9.215 126.445 9.785 ;
  END
 END i22
 PIN i23
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 10.735 126.445 11.305 ;
  END
 END i23
 PIN i24
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 11.495 126.445 12.065 ;
  END
 END i24
 PIN i25
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 12.255 126.445 12.825 ;
  END
 END i25
 PIN i26
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 13.015 126.445 13.585 ;
  END
 END i26
 PIN i27
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 8.075 125.685 8.645 ;
  END
 END i27
 PIN i28
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 7.695 126.445 8.265 ;
  END
 END i28
 PIN i29
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 7.315 125.685 7.885 ;
  END
 END i29
 PIN i30
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 6.935 126.445 7.505 ;
  END
 END i30
 PIN i31
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 6.555 125.685 7.125 ;
  END
 END i31
 PIN i32
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 13.775 126.445 14.345 ;
  END
 END i32
 PIN i33
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 15.295 126.445 15.865 ;
  END
 END i33
 PIN i34
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 16.055 126.445 16.625 ;
  END
 END i34
 PIN i35
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 16.815 126.445 17.385 ;
  END
 END i35
 OBS
  LAYER metal1 ;
   RECT 0 0 129.58 70.11 ;
  LAYER via1 ;
   RECT 0 0 129.58 70.11 ;
  LAYER metal2 ;
   RECT 0 0 129.58 70.11 ;
  LAYER via2 ;
   RECT 0 0 129.58 70.11 ;
  LAYER metal3 ;
   RECT 0 0 129.58 70.11 ;
  LAYER via3 ;
   RECT 0 0 129.58 70.11 ;
  LAYER metal4 ;
   RECT 0 0 129.58 70.11 ;
 END
END block_341x369_82

MACRO block_414x1746_310
 CLASS BLOCK ;
 FOREIGN block_414x1746_310 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 157.32 BY 331.74 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 326.515 131.005 327.085 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 322.335 131.005 322.905 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 285.665 131.005 286.235 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 281.485 131.005 282.055 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 277.495 131.005 278.065 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 273.315 131.005 273.885 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 269.325 131.005 269.895 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 265.145 131.005 265.715 ;
  END
 END o7
 PIN o8
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 261.155 131.005 261.725 ;
  END
 END o8
 PIN o9
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 238.735 131.005 239.305 ;
  END
 END o9
 PIN o10
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 234.745 131.005 235.315 ;
  END
 END o10
 PIN o11
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 230.565 131.005 231.135 ;
  END
 END o11
 PIN o12
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 318.345 131.005 318.915 ;
  END
 END o12
 PIN o13
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 226.575 131.005 227.145 ;
  END
 END o13
 PIN o14
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 222.395 131.005 222.965 ;
  END
 END o14
 PIN o15
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 218.405 131.005 218.975 ;
  END
 END o15
 PIN o16
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 214.225 131.005 214.795 ;
  END
 END o16
 PIN o17
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 210.235 131.005 210.805 ;
  END
 END o17
 PIN o18
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 206.055 131.005 206.625 ;
  END
 END o18
 PIN o19
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 202.065 131.005 202.635 ;
  END
 END o19
 PIN o20
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 197.885 131.005 198.455 ;
  END
 END o20
 PIN o21
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 193.895 131.005 194.465 ;
  END
 END o21
 PIN o22
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 189.715 131.005 190.285 ;
  END
 END o22
 PIN o23
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 314.165 131.005 314.735 ;
  END
 END o23
 PIN o24
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 185.725 131.005 186.295 ;
  END
 END o24
 PIN o25
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 181.545 131.005 182.115 ;
  END
 END o25
 PIN o26
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 177.555 131.005 178.125 ;
  END
 END o26
 PIN o27
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 149.245 131.005 149.815 ;
  END
 END o27
 PIN o28
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 145.255 131.005 145.825 ;
  END
 END o28
 PIN o29
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 141.075 131.005 141.645 ;
  END
 END o29
 PIN o30
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 137.085 131.005 137.655 ;
  END
 END o30
 PIN o31
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 132.905 131.005 133.475 ;
  END
 END o31
 PIN o32
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 128.915 131.005 129.485 ;
  END
 END o32
 PIN o33
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 124.735 131.005 125.305 ;
  END
 END o33
 PIN o34
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 310.175 131.005 310.745 ;
  END
 END o34
 PIN o35
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 120.745 131.005 121.315 ;
  END
 END o35
 PIN o36
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 116.565 131.005 117.135 ;
  END
 END o36
 PIN o37
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 112.575 131.005 113.145 ;
  END
 END o37
 PIN o38
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 108.395 131.005 108.965 ;
  END
 END o38
 PIN o39
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 104.405 131.005 104.975 ;
  END
 END o39
 PIN o40
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 100.225 131.005 100.795 ;
  END
 END o40
 PIN o41
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 96.235 131.005 96.805 ;
  END
 END o41
 PIN o42
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 92.055 131.005 92.625 ;
  END
 END o42
 PIN o43
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 88.065 131.005 88.635 ;
  END
 END o43
 PIN o44
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 65.645 131.005 66.215 ;
  END
 END o44
 PIN o45
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 305.995 131.005 306.565 ;
  END
 END o45
 PIN o46
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 61.655 131.005 62.225 ;
  END
 END o46
 PIN o47
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 57.475 131.005 58.045 ;
  END
 END o47
 PIN o48
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 53.485 131.005 54.055 ;
  END
 END o48
 PIN o49
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 49.305 131.005 49.875 ;
  END
 END o49
 PIN o50
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 45.315 131.005 45.885 ;
  END
 END o50
 PIN o51
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 41.135 131.005 41.705 ;
  END
 END o51
 PIN o52
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 37.145 131.005 37.715 ;
  END
 END o52
 PIN o53
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 32.965 131.005 33.535 ;
  END
 END o53
 PIN o54
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 28.975 131.005 29.545 ;
  END
 END o54
 PIN o55
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 24.795 131.005 25.365 ;
  END
 END o55
 PIN o56
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 302.005 131.005 302.575 ;
  END
 END o56
 PIN o57
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 20.805 131.005 21.375 ;
  END
 END o57
 PIN o58
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 16.625 131.005 17.195 ;
  END
 END o58
 PIN o59
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 12.635 131.005 13.205 ;
  END
 END o59
 PIN o60
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 8.455 131.005 9.025 ;
  END
 END o60
 PIN o61
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 4.465 131.005 5.035 ;
  END
 END o61
 PIN o62
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 297.825 131.005 298.395 ;
  END
 END o62
 PIN o63
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 293.835 131.005 294.405 ;
  END
 END o63
 PIN o64
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 289.655 131.005 290.225 ;
  END
 END o64
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 153.615 174.515 154.185 175.085 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 153.615 157.415 154.185 157.985 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 153.615 169.195 154.185 169.765 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 152.855 174.135 153.425 174.705 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 152.855 174.895 153.425 175.465 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 153.615 175.275 154.185 175.845 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 153.615 165.585 154.185 166.155 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 153.615 152.475 154.185 153.045 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 153.615 158.175 154.185 158.745 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 153.615 156.085 154.185 156.655 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 153.615 153.615 154.185 154.185 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 152.855 152.095 153.425 152.665 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 143.735 175.655 144.305 176.225 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 143.735 162.355 144.305 162.925 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 328.225 131.005 328.795 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 324.045 131.005 324.615 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 287.375 131.005 287.945 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 283.195 131.005 283.765 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 279.205 131.005 279.775 ;
  END
 END i18
 PIN i19
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 275.025 131.005 275.595 ;
  END
 END i19
 PIN i20
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 271.035 131.005 271.605 ;
  END
 END i20
 PIN i21
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 266.855 131.005 267.425 ;
  END
 END i21
 PIN i22
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 262.865 131.005 263.435 ;
  END
 END i22
 PIN i23
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 240.445 131.005 241.015 ;
  END
 END i23
 PIN i24
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 236.455 131.005 237.025 ;
  END
 END i24
 PIN i25
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 232.275 131.005 232.845 ;
  END
 END i25
 PIN i26
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 320.055 131.005 320.625 ;
  END
 END i26
 PIN i27
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 228.285 131.005 228.855 ;
  END
 END i27
 PIN i28
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 224.105 131.005 224.675 ;
  END
 END i28
 PIN i29
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 220.115 131.005 220.685 ;
  END
 END i29
 PIN i30
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 215.935 131.005 216.505 ;
  END
 END i30
 PIN i31
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 211.945 131.005 212.515 ;
  END
 END i31
 PIN i32
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 207.765 131.005 208.335 ;
  END
 END i32
 PIN i33
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 203.775 131.005 204.345 ;
  END
 END i33
 PIN i34
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 199.595 131.005 200.165 ;
  END
 END i34
 PIN i35
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 195.605 131.005 196.175 ;
  END
 END i35
 PIN i36
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 191.425 131.005 191.995 ;
  END
 END i36
 PIN i37
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 315.875 131.005 316.445 ;
  END
 END i37
 PIN i38
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 187.435 131.005 188.005 ;
  END
 END i38
 PIN i39
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 183.255 131.005 183.825 ;
  END
 END i39
 PIN i40
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 179.265 131.005 179.835 ;
  END
 END i40
 PIN i41
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 147.535 131.005 148.105 ;
  END
 END i41
 PIN i42
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 143.545 131.005 144.115 ;
  END
 END i42
 PIN i43
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 139.365 131.005 139.935 ;
  END
 END i43
 PIN i44
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 135.375 131.005 135.945 ;
  END
 END i44
 PIN i45
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 131.195 131.005 131.765 ;
  END
 END i45
 PIN i46
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 127.205 131.005 127.775 ;
  END
 END i46
 PIN i47
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 123.025 131.005 123.595 ;
  END
 END i47
 PIN i48
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 311.885 131.005 312.455 ;
  END
 END i48
 PIN i49
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 119.035 131.005 119.605 ;
  END
 END i49
 PIN i50
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 114.855 131.005 115.425 ;
  END
 END i50
 PIN i51
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 110.865 131.005 111.435 ;
  END
 END i51
 PIN i52
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 106.685 131.005 107.255 ;
  END
 END i52
 PIN i53
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 102.695 131.005 103.265 ;
  END
 END i53
 PIN i54
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 98.515 131.005 99.085 ;
  END
 END i54
 PIN i55
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 94.525 131.005 95.095 ;
  END
 END i55
 PIN i56
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 90.345 131.005 90.915 ;
  END
 END i56
 PIN i57
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 86.355 131.005 86.925 ;
  END
 END i57
 PIN i58
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 63.935 131.005 64.505 ;
  END
 END i58
 PIN i59
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 307.705 131.005 308.275 ;
  END
 END i59
 PIN i60
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 59.945 131.005 60.515 ;
  END
 END i60
 PIN i61
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 55.765 131.005 56.335 ;
  END
 END i61
 PIN i62
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 51.775 131.005 52.345 ;
  END
 END i62
 PIN i63
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 47.595 131.005 48.165 ;
  END
 END i63
 PIN i64
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 43.605 131.005 44.175 ;
  END
 END i64
 PIN i65
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 39.425 131.005 39.995 ;
  END
 END i65
 PIN i66
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 35.435 131.005 36.005 ;
  END
 END i66
 PIN i67
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 31.255 131.005 31.825 ;
  END
 END i67
 PIN i68
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 27.265 131.005 27.835 ;
  END
 END i68
 PIN i69
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 23.085 131.005 23.655 ;
  END
 END i69
 PIN i70
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 303.715 131.005 304.285 ;
  END
 END i70
 PIN i71
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 19.095 131.005 19.665 ;
  END
 END i71
 PIN i72
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 14.915 131.005 15.485 ;
  END
 END i72
 PIN i73
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 10.925 131.005 11.495 ;
  END
 END i73
 PIN i74
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 6.745 131.005 7.315 ;
  END
 END i74
 PIN i75
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 2.755 131.005 3.325 ;
  END
 END i75
 PIN i76
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 299.535 131.005 300.105 ;
  END
 END i76
 PIN i77
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 295.545 131.005 296.115 ;
  END
 END i77
 PIN i78
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.435 291.365 131.005 291.935 ;
  END
 END i78
 PIN i79
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 285.095 130.245 285.665 ;
  END
 END i79
 PIN i80
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 280.915 130.245 281.485 ;
  END
 END i80
 PIN i81
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 276.925 130.245 277.495 ;
  END
 END i81
 PIN i82
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 297.255 130.245 297.825 ;
  END
 END i82
 PIN i83
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 293.265 130.245 293.835 ;
  END
 END i83
 PIN i84
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 217.835 130.245 218.405 ;
  END
 END i84
 PIN i85
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 213.655 130.245 214.225 ;
  END
 END i85
 PIN i86
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 209.665 130.245 210.235 ;
  END
 END i86
 PIN i87
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 205.485 130.245 206.055 ;
  END
 END i87
 PIN i88
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 226.005 130.245 226.575 ;
  END
 END i88
 PIN i89
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 108.965 130.245 109.535 ;
  END
 END i89
 PIN i90
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 113.145 130.245 113.715 ;
  END
 END i90
 PIN i91
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 117.135 130.245 117.705 ;
  END
 END i91
 PIN i92
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 121.315 130.245 121.885 ;
  END
 END i92
 PIN i93
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 100.795 130.245 101.365 ;
  END
 END i93
 PIN i94
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 41.705 130.245 42.275 ;
  END
 END i94
 PIN i95
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 45.885 130.245 46.455 ;
  END
 END i95
 PIN i96
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 49.875 130.245 50.445 ;
  END
 END i96
 PIN i97
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 33.535 130.245 34.105 ;
  END
 END i97
 PIN i98
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 54.055 130.245 54.625 ;
  END
 END i98
 PIN i99
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 289.085 130.245 289.655 ;
  END
 END i99
 PIN i100
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 221.825 130.245 222.395 ;
  END
 END i100
 PIN i101
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 104.975 130.245 105.545 ;
  END
 END i101
 PIN i102
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 37.715 130.245 38.285 ;
  END
 END i102
 PIN i103
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 138.795 175.655 139.365 176.225 ;
  END
 END i103
 PIN i104
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 138.795 162.355 139.365 162.925 ;
  END
 END i104
 PIN i105
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 327.655 130.245 328.225 ;
  END
 END i105
 PIN i106
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 323.475 130.245 324.045 ;
  END
 END i106
 PIN i107
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 286.805 130.245 287.375 ;
  END
 END i107
 PIN i108
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 282.625 130.245 283.195 ;
  END
 END i108
 PIN i109
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 278.635 130.245 279.205 ;
  END
 END i109
 PIN i110
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 274.455 130.245 275.025 ;
  END
 END i110
 PIN i111
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 270.465 130.245 271.035 ;
  END
 END i111
 PIN i112
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 266.285 130.245 266.855 ;
  END
 END i112
 PIN i113
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 262.295 130.245 262.865 ;
  END
 END i113
 PIN i114
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 239.875 130.245 240.445 ;
  END
 END i114
 PIN i115
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 235.885 130.245 236.455 ;
  END
 END i115
 PIN i116
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 231.705 130.245 232.275 ;
  END
 END i116
 PIN i117
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 319.485 130.245 320.055 ;
  END
 END i117
 PIN i118
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 227.715 130.245 228.285 ;
  END
 END i118
 PIN i119
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 223.535 130.245 224.105 ;
  END
 END i119
 PIN i120
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 219.545 130.245 220.115 ;
  END
 END i120
 PIN i121
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 215.365 130.245 215.935 ;
  END
 END i121
 PIN i122
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 211.375 130.245 211.945 ;
  END
 END i122
 PIN i123
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 207.195 130.245 207.765 ;
  END
 END i123
 PIN i124
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 203.205 130.245 203.775 ;
  END
 END i124
 PIN i125
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 199.025 130.245 199.595 ;
  END
 END i125
 PIN i126
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 195.035 130.245 195.605 ;
  END
 END i126
 PIN i127
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 190.855 130.245 191.425 ;
  END
 END i127
 PIN i128
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 315.305 130.245 315.875 ;
  END
 END i128
 PIN i129
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 186.865 130.245 187.435 ;
  END
 END i129
 PIN i130
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 182.685 130.245 183.255 ;
  END
 END i130
 PIN i131
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 178.695 130.245 179.265 ;
  END
 END i131
 PIN i132
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 148.105 130.245 148.675 ;
  END
 END i132
 PIN i133
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 144.115 130.245 144.685 ;
  END
 END i133
 PIN i134
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 139.935 130.245 140.505 ;
  END
 END i134
 PIN i135
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 135.945 130.245 136.515 ;
  END
 END i135
 PIN i136
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 131.765 130.245 132.335 ;
  END
 END i136
 PIN i137
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 127.775 130.245 128.345 ;
  END
 END i137
 PIN i138
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 123.595 130.245 124.165 ;
  END
 END i138
 PIN i139
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 311.315 130.245 311.885 ;
  END
 END i139
 PIN i140
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 119.605 130.245 120.175 ;
  END
 END i140
 PIN i141
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 115.425 130.245 115.995 ;
  END
 END i141
 PIN i142
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 111.435 130.245 112.005 ;
  END
 END i142
 PIN i143
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 107.255 130.245 107.825 ;
  END
 END i143
 PIN i144
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 103.265 130.245 103.835 ;
  END
 END i144
 PIN i145
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 99.085 130.245 99.655 ;
  END
 END i145
 PIN i146
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 95.095 130.245 95.665 ;
  END
 END i146
 PIN i147
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 90.915 130.245 91.485 ;
  END
 END i147
 PIN i148
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 86.925 130.245 87.495 ;
  END
 END i148
 PIN i149
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 64.505 130.245 65.075 ;
  END
 END i149
 PIN i150
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 307.135 130.245 307.705 ;
  END
 END i150
 PIN i151
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 60.515 130.245 61.085 ;
  END
 END i151
 PIN i152
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 56.335 130.245 56.905 ;
  END
 END i152
 PIN i153
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 52.345 130.245 52.915 ;
  END
 END i153
 PIN i154
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 48.165 130.245 48.735 ;
  END
 END i154
 PIN i155
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 44.175 130.245 44.745 ;
  END
 END i155
 PIN i156
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 39.995 130.245 40.565 ;
  END
 END i156
 PIN i157
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 36.005 130.245 36.575 ;
  END
 END i157
 PIN i158
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 31.825 130.245 32.395 ;
  END
 END i158
 PIN i159
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 27.835 130.245 28.405 ;
  END
 END i159
 PIN i160
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 23.655 130.245 24.225 ;
  END
 END i160
 PIN i161
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 303.145 130.245 303.715 ;
  END
 END i161
 PIN i162
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 19.665 130.245 20.235 ;
  END
 END i162
 PIN i163
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 15.485 130.245 16.055 ;
  END
 END i163
 PIN i164
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 11.495 130.245 12.065 ;
  END
 END i164
 PIN i165
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 7.315 130.245 7.885 ;
  END
 END i165
 PIN i166
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 3.325 130.245 3.895 ;
  END
 END i166
 PIN i167
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 298.965 130.245 299.535 ;
  END
 END i167
 PIN i168
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 294.975 130.245 295.545 ;
  END
 END i168
 PIN i169
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 290.795 130.245 291.365 ;
  END
 END i169
 PIN i170
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 153.615 168.055 154.185 168.625 ;
  END
 END i170
 PIN i171
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 152.855 167.675 153.425 168.245 ;
  END
 END i171
 PIN i172
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 327.085 129.485 327.655 ;
  END
 END i172
 PIN i173
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 322.905 129.485 323.475 ;
  END
 END i173
 PIN i174
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 286.235 129.485 286.805 ;
  END
 END i174
 PIN i175
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 282.055 129.485 282.625 ;
  END
 END i175
 PIN i176
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 278.065 129.485 278.635 ;
  END
 END i176
 PIN i177
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 273.885 129.485 274.455 ;
  END
 END i177
 PIN i178
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 269.895 129.485 270.465 ;
  END
 END i178
 PIN i179
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 265.715 129.485 266.285 ;
  END
 END i179
 PIN i180
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 261.725 129.485 262.295 ;
  END
 END i180
 PIN i181
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 239.305 129.485 239.875 ;
  END
 END i181
 PIN i182
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 235.315 129.485 235.885 ;
  END
 END i182
 PIN i183
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 231.135 129.485 231.705 ;
  END
 END i183
 PIN i184
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 318.915 129.485 319.485 ;
  END
 END i184
 PIN i185
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 227.145 129.485 227.715 ;
  END
 END i185
 PIN i186
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 222.965 129.485 223.535 ;
  END
 END i186
 PIN i187
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 218.975 129.485 219.545 ;
  END
 END i187
 PIN i188
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 214.795 129.485 215.365 ;
  END
 END i188
 PIN i189
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 210.805 129.485 211.375 ;
  END
 END i189
 PIN i190
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 206.625 129.485 207.195 ;
  END
 END i190
 PIN i191
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 202.635 129.485 203.205 ;
  END
 END i191
 PIN i192
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 198.455 129.485 199.025 ;
  END
 END i192
 PIN i193
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 194.465 129.485 195.035 ;
  END
 END i193
 PIN i194
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 190.285 129.485 190.855 ;
  END
 END i194
 PIN i195
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 314.735 129.485 315.305 ;
  END
 END i195
 PIN i196
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 186.295 129.485 186.865 ;
  END
 END i196
 PIN i197
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 182.115 129.485 182.685 ;
  END
 END i197
 PIN i198
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 178.125 129.485 178.695 ;
  END
 END i198
 PIN i199
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 148.675 129.485 149.245 ;
  END
 END i199
 PIN i200
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 144.685 129.485 145.255 ;
  END
 END i200
 PIN i201
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 140.505 129.485 141.075 ;
  END
 END i201
 PIN i202
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 136.515 129.485 137.085 ;
  END
 END i202
 PIN i203
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 132.335 129.485 132.905 ;
  END
 END i203
 PIN i204
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 128.345 129.485 128.915 ;
  END
 END i204
 PIN i205
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 124.165 129.485 124.735 ;
  END
 END i205
 PIN i206
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 310.745 129.485 311.315 ;
  END
 END i206
 PIN i207
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 120.175 129.485 120.745 ;
  END
 END i207
 PIN i208
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 115.995 129.485 116.565 ;
  END
 END i208
 PIN i209
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 112.005 129.485 112.575 ;
  END
 END i209
 PIN i210
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 107.825 129.485 108.395 ;
  END
 END i210
 PIN i211
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 103.835 129.485 104.405 ;
  END
 END i211
 PIN i212
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 99.655 129.485 100.225 ;
  END
 END i212
 PIN i213
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 95.665 129.485 96.235 ;
  END
 END i213
 PIN i214
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 91.485 129.485 92.055 ;
  END
 END i214
 PIN i215
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 87.495 129.485 88.065 ;
  END
 END i215
 PIN i216
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 65.075 129.485 65.645 ;
  END
 END i216
 PIN i217
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 306.565 129.485 307.135 ;
  END
 END i217
 PIN i218
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 61.085 129.485 61.655 ;
  END
 END i218
 PIN i219
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 56.905 129.485 57.475 ;
  END
 END i219
 PIN i220
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 52.915 129.485 53.485 ;
  END
 END i220
 PIN i221
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 48.735 129.485 49.305 ;
  END
 END i221
 PIN i222
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 44.745 129.485 45.315 ;
  END
 END i222
 PIN i223
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 40.565 129.485 41.135 ;
  END
 END i223
 PIN i224
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 36.575 129.485 37.145 ;
  END
 END i224
 PIN i225
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 32.395 129.485 32.965 ;
  END
 END i225
 PIN i226
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 28.405 129.485 28.975 ;
  END
 END i226
 PIN i227
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 24.225 129.485 24.795 ;
  END
 END i227
 PIN i228
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 302.575 129.485 303.145 ;
  END
 END i228
 PIN i229
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 20.235 129.485 20.805 ;
  END
 END i229
 PIN i230
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 16.055 129.485 16.625 ;
  END
 END i230
 PIN i231
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 12.065 129.485 12.635 ;
  END
 END i231
 PIN i232
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 7.885 129.485 8.455 ;
  END
 END i232
 PIN i233
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 3.895 129.485 4.465 ;
  END
 END i233
 PIN i234
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 298.395 129.485 298.965 ;
  END
 END i234
 PIN i235
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 294.405 129.485 294.975 ;
  END
 END i235
 PIN i236
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 290.225 129.485 290.795 ;
  END
 END i236
 PIN i237
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 152.475 175.655 153.045 176.225 ;
  END
 END i237
 PIN i238
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 151.335 175.655 151.905 176.225 ;
  END
 END i238
 PIN i239
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 149.815 175.655 150.385 176.225 ;
  END
 END i239
 PIN i240
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 147.915 175.655 148.485 176.225 ;
  END
 END i240
 PIN i241
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 152.475 162.355 153.045 162.925 ;
  END
 END i241
 PIN i242
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 151.335 162.355 151.905 162.925 ;
  END
 END i242
 PIN i243
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 149.815 162.355 150.385 162.925 ;
  END
 END i243
 PIN i244
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 147.915 162.355 148.485 162.925 ;
  END
 END i244
 OBS
  LAYER metal1 ;
   RECT 0.0 0.0 134.14 1.71 ;
   RECT 0.0 1.71 134.14 3.42 ;
   RECT 0.0 3.42 134.14 5.13 ;
   RECT 0.0 5.13 134.14 6.84 ;
   RECT 0.0 6.84 134.14 8.55 ;
   RECT 0.0 8.55 134.14 10.26 ;
   RECT 0.0 10.26 134.14 11.97 ;
   RECT 0.0 11.97 134.14 13.68 ;
   RECT 0.0 13.68 134.14 15.39 ;
   RECT 0.0 15.39 134.14 17.1 ;
   RECT 0.0 17.1 134.14 18.81 ;
   RECT 0.0 18.81 134.14 20.52 ;
   RECT 0.0 20.52 134.14 22.23 ;
   RECT 0.0 22.23 134.14 23.94 ;
   RECT 0.0 23.94 134.14 25.65 ;
   RECT 0.0 25.65 134.14 27.36 ;
   RECT 0.0 27.36 134.14 29.07 ;
   RECT 0.0 29.07 134.14 30.78 ;
   RECT 0.0 30.78 134.14 32.49 ;
   RECT 0.0 32.49 134.14 34.2 ;
   RECT 0.0 34.2 134.14 35.91 ;
   RECT 0.0 35.91 134.14 37.62 ;
   RECT 0.0 37.62 134.14 39.33 ;
   RECT 0.0 39.33 134.14 41.04 ;
   RECT 0.0 41.04 134.14 42.75 ;
   RECT 0.0 42.75 134.14 44.46 ;
   RECT 0.0 44.46 134.14 46.17 ;
   RECT 0.0 46.17 134.14 47.88 ;
   RECT 0.0 47.88 134.14 49.59 ;
   RECT 0.0 49.59 134.14 51.3 ;
   RECT 0.0 51.3 134.14 53.01 ;
   RECT 0.0 53.01 134.14 54.72 ;
   RECT 0.0 54.72 134.14 56.43 ;
   RECT 0.0 56.43 134.14 58.14 ;
   RECT 0.0 58.14 134.14 59.85 ;
   RECT 0.0 59.85 134.14 61.56 ;
   RECT 0.0 61.56 134.14 63.27 ;
   RECT 0.0 63.27 134.14 64.98 ;
   RECT 0.0 64.98 134.14 66.69 ;
   RECT 0.0 66.69 134.14 68.4 ;
   RECT 0.0 68.4 134.14 70.11 ;
   RECT 0.0 70.11 134.14 71.82 ;
   RECT 0.0 71.82 134.14 73.53 ;
   RECT 0.0 73.53 134.14 75.24 ;
   RECT 0.0 75.24 134.14 76.95 ;
   RECT 0.0 76.95 134.14 78.66 ;
   RECT 0.0 78.66 134.14 80.37 ;
   RECT 0.0 80.37 134.14 82.08 ;
   RECT 0.0 82.08 134.14 83.79 ;
   RECT 0.0 83.79 134.14 85.5 ;
   RECT 0.0 85.5 134.14 87.21 ;
   RECT 0.0 87.21 134.14 88.92 ;
   RECT 0.0 88.92 134.14 90.63 ;
   RECT 0.0 90.63 134.14 92.34 ;
   RECT 0.0 92.34 134.14 94.05 ;
   RECT 0.0 94.05 134.14 95.76 ;
   RECT 0.0 95.76 134.14 97.47 ;
   RECT 0.0 97.47 134.14 99.18 ;
   RECT 0.0 99.18 134.14 100.89 ;
   RECT 0.0 100.89 134.14 102.6 ;
   RECT 0.0 102.6 134.14 104.31 ;
   RECT 0.0 104.31 134.14 106.02 ;
   RECT 0.0 106.02 134.14 107.73 ;
   RECT 0.0 107.73 134.14 109.44 ;
   RECT 0.0 109.44 134.14 111.15 ;
   RECT 0.0 111.15 134.14 112.86 ;
   RECT 0.0 112.86 134.14 114.57 ;
   RECT 0.0 114.57 134.14 116.28 ;
   RECT 0.0 116.28 134.14 117.99 ;
   RECT 0.0 117.99 134.14 119.7 ;
   RECT 0.0 119.7 134.14 121.41 ;
   RECT 0.0 121.41 134.14 123.12 ;
   RECT 0.0 123.12 134.14 124.83 ;
   RECT 0.0 124.83 134.14 126.54 ;
   RECT 0.0 126.54 134.14 128.25 ;
   RECT 0.0 128.25 134.14 129.96 ;
   RECT 0.0 129.96 134.14 131.67 ;
   RECT 0.0 131.67 134.14 133.38 ;
   RECT 0.0 133.38 134.14 135.09 ;
   RECT 0.0 135.09 134.14 136.8 ;
   RECT 0.0 136.8 134.14 138.51 ;
   RECT 0.0 138.51 134.14 140.22 ;
   RECT 0.0 140.22 134.14 141.93 ;
   RECT 0.0 141.93 134.14 143.64 ;
   RECT 0.0 143.64 134.14 145.35 ;
   RECT 0.0 145.35 134.14 147.06 ;
   RECT 0.0 147.06 134.14 148.77 ;
   RECT 0.0 148.77 157.32 150.48 ;
   RECT 0.0 150.48 157.32 152.19 ;
   RECT 0.0 152.19 157.32 153.9 ;
   RECT 0.0 153.9 157.32 155.61 ;
   RECT 0.0 155.61 157.32 157.32 ;
   RECT 0.0 157.32 157.32 159.03 ;
   RECT 0.0 159.03 157.32 160.74 ;
   RECT 0.0 160.74 157.32 162.45 ;
   RECT 0.0 162.45 157.32 164.16 ;
   RECT 0.0 164.16 157.32 165.87 ;
   RECT 0.0 165.87 157.32 167.58 ;
   RECT 0.0 167.58 157.32 169.29 ;
   RECT 0.0 169.29 157.32 171.0 ;
   RECT 0.0 171.0 157.32 172.71 ;
   RECT 0.0 172.71 157.32 174.42 ;
   RECT 0.0 174.42 157.32 176.13 ;
   RECT 0.0 176.13 157.32 177.84 ;
   RECT 0.0 177.84 134.14 179.55 ;
   RECT 0.0 179.55 134.14 181.26 ;
   RECT 0.0 181.26 134.14 182.97 ;
   RECT 0.0 182.97 134.14 184.68 ;
   RECT 0.0 184.68 134.14 186.39 ;
   RECT 0.0 186.39 134.14 188.1 ;
   RECT 0.0 188.1 134.14 189.81 ;
   RECT 0.0 189.81 134.14 191.52 ;
   RECT 0.0 191.52 134.14 193.23 ;
   RECT 0.0 193.23 134.14 194.94 ;
   RECT 0.0 194.94 134.14 196.65 ;
   RECT 0.0 196.65 134.14 198.36 ;
   RECT 0.0 198.36 134.14 200.07 ;
   RECT 0.0 200.07 134.14 201.78 ;
   RECT 0.0 201.78 134.14 203.49 ;
   RECT 0.0 203.49 134.14 205.2 ;
   RECT 0.0 205.2 134.14 206.91 ;
   RECT 0.0 206.91 134.14 208.62 ;
   RECT 0.0 208.62 134.14 210.33 ;
   RECT 0.0 210.33 134.14 212.04 ;
   RECT 0.0 212.04 134.14 213.75 ;
   RECT 0.0 213.75 134.14 215.46 ;
   RECT 0.0 215.46 134.14 217.17 ;
   RECT 0.0 217.17 134.14 218.88 ;
   RECT 0.0 218.88 134.14 220.59 ;
   RECT 0.0 220.59 134.14 222.3 ;
   RECT 0.0 222.3 134.14 224.01 ;
   RECT 0.0 224.01 134.14 225.72 ;
   RECT 0.0 225.72 134.14 227.43 ;
   RECT 0.0 227.43 134.14 229.14 ;
   RECT 0.0 229.14 134.14 230.85 ;
   RECT 0.0 230.85 134.14 232.56 ;
   RECT 0.0 232.56 134.14 234.27 ;
   RECT 0.0 234.27 134.14 235.98 ;
   RECT 0.0 235.98 134.14 237.69 ;
   RECT 0.0 237.69 134.14 239.4 ;
   RECT 0.0 239.4 134.14 241.11 ;
   RECT 0.0 241.11 134.14 242.82 ;
   RECT 0.0 242.82 134.14 244.53 ;
   RECT 0.0 244.53 134.14 246.24 ;
   RECT 0.0 246.24 134.14 247.95 ;
   RECT 0.0 247.95 134.14 249.66 ;
   RECT 0.0 249.66 134.14 251.37 ;
   RECT 0.0 251.37 134.14 253.08 ;
   RECT 0.0 253.08 134.14 254.79 ;
   RECT 0.0 254.79 134.14 256.5 ;
   RECT 0.0 256.5 134.14 258.21 ;
   RECT 0.0 258.21 134.14 259.92 ;
   RECT 0.0 259.92 134.14 261.63 ;
   RECT 0.0 261.63 134.14 263.34 ;
   RECT 0.0 263.34 134.14 265.05 ;
   RECT 0.0 265.05 134.14 266.76 ;
   RECT 0.0 266.76 134.14 268.47 ;
   RECT 0.0 268.47 134.14 270.18 ;
   RECT 0.0 270.18 134.14 271.89 ;
   RECT 0.0 271.89 134.14 273.6 ;
   RECT 0.0 273.6 134.14 275.31 ;
   RECT 0.0 275.31 134.14 277.02 ;
   RECT 0.0 277.02 134.14 278.73 ;
   RECT 0.0 278.73 134.14 280.44 ;
   RECT 0.0 280.44 134.14 282.15 ;
   RECT 0.0 282.15 134.14 283.86 ;
   RECT 0.0 283.86 134.14 285.57 ;
   RECT 0.0 285.57 134.14 287.28 ;
   RECT 0.0 287.28 134.14 288.99 ;
   RECT 0.0 288.99 134.14 290.7 ;
   RECT 0.0 290.7 134.14 292.41 ;
   RECT 0.0 292.41 134.14 294.12 ;
   RECT 0.0 294.12 134.14 295.83 ;
   RECT 0.0 295.83 134.14 297.54 ;
   RECT 0.0 297.54 134.14 299.25 ;
   RECT 0.0 299.25 134.14 300.96 ;
   RECT 0.0 300.96 134.14 302.67 ;
   RECT 0.0 302.67 134.14 304.38 ;
   RECT 0.0 304.38 134.14 306.09 ;
   RECT 0.0 306.09 134.14 307.8 ;
   RECT 0.0 307.8 134.14 309.51 ;
   RECT 0.0 309.51 134.14 311.22 ;
   RECT 0.0 311.22 134.14 312.93 ;
   RECT 0.0 312.93 134.14 314.64 ;
   RECT 0.0 314.64 134.14 316.35 ;
   RECT 0.0 316.35 134.14 318.06 ;
   RECT 0.0 318.06 134.14 319.77 ;
   RECT 0.0 319.77 134.14 321.48 ;
   RECT 0.0 321.48 134.14 323.19 ;
   RECT 0.0 323.19 134.14 324.9 ;
   RECT 0.0 324.9 134.14 326.61 ;
   RECT 0.0 326.61 134.14 328.32 ;
   RECT 0.0 328.32 134.14 330.03 ;
   RECT 0.0 330.03 134.14 331.74 ;
  LAYER via1 ;
   RECT 0.0 0.0 134.14 1.71 ;
   RECT 0.0 1.71 134.14 3.42 ;
   RECT 0.0 3.42 134.14 5.13 ;
   RECT 0.0 5.13 134.14 6.84 ;
   RECT 0.0 6.84 134.14 8.55 ;
   RECT 0.0 8.55 134.14 10.26 ;
   RECT 0.0 10.26 134.14 11.97 ;
   RECT 0.0 11.97 134.14 13.68 ;
   RECT 0.0 13.68 134.14 15.39 ;
   RECT 0.0 15.39 134.14 17.1 ;
   RECT 0.0 17.1 134.14 18.81 ;
   RECT 0.0 18.81 134.14 20.52 ;
   RECT 0.0 20.52 134.14 22.23 ;
   RECT 0.0 22.23 134.14 23.94 ;
   RECT 0.0 23.94 134.14 25.65 ;
   RECT 0.0 25.65 134.14 27.36 ;
   RECT 0.0 27.36 134.14 29.07 ;
   RECT 0.0 29.07 134.14 30.78 ;
   RECT 0.0 30.78 134.14 32.49 ;
   RECT 0.0 32.49 134.14 34.2 ;
   RECT 0.0 34.2 134.14 35.91 ;
   RECT 0.0 35.91 134.14 37.62 ;
   RECT 0.0 37.62 134.14 39.33 ;
   RECT 0.0 39.33 134.14 41.04 ;
   RECT 0.0 41.04 134.14 42.75 ;
   RECT 0.0 42.75 134.14 44.46 ;
   RECT 0.0 44.46 134.14 46.17 ;
   RECT 0.0 46.17 134.14 47.88 ;
   RECT 0.0 47.88 134.14 49.59 ;
   RECT 0.0 49.59 134.14 51.3 ;
   RECT 0.0 51.3 134.14 53.01 ;
   RECT 0.0 53.01 134.14 54.72 ;
   RECT 0.0 54.72 134.14 56.43 ;
   RECT 0.0 56.43 134.14 58.14 ;
   RECT 0.0 58.14 134.14 59.85 ;
   RECT 0.0 59.85 134.14 61.56 ;
   RECT 0.0 61.56 134.14 63.27 ;
   RECT 0.0 63.27 134.14 64.98 ;
   RECT 0.0 64.98 134.14 66.69 ;
   RECT 0.0 66.69 134.14 68.4 ;
   RECT 0.0 68.4 134.14 70.11 ;
   RECT 0.0 70.11 134.14 71.82 ;
   RECT 0.0 71.82 134.14 73.53 ;
   RECT 0.0 73.53 134.14 75.24 ;
   RECT 0.0 75.24 134.14 76.95 ;
   RECT 0.0 76.95 134.14 78.66 ;
   RECT 0.0 78.66 134.14 80.37 ;
   RECT 0.0 80.37 134.14 82.08 ;
   RECT 0.0 82.08 134.14 83.79 ;
   RECT 0.0 83.79 134.14 85.5 ;
   RECT 0.0 85.5 134.14 87.21 ;
   RECT 0.0 87.21 134.14 88.92 ;
   RECT 0.0 88.92 134.14 90.63 ;
   RECT 0.0 90.63 134.14 92.34 ;
   RECT 0.0 92.34 134.14 94.05 ;
   RECT 0.0 94.05 134.14 95.76 ;
   RECT 0.0 95.76 134.14 97.47 ;
   RECT 0.0 97.47 134.14 99.18 ;
   RECT 0.0 99.18 134.14 100.89 ;
   RECT 0.0 100.89 134.14 102.6 ;
   RECT 0.0 102.6 134.14 104.31 ;
   RECT 0.0 104.31 134.14 106.02 ;
   RECT 0.0 106.02 134.14 107.73 ;
   RECT 0.0 107.73 134.14 109.44 ;
   RECT 0.0 109.44 134.14 111.15 ;
   RECT 0.0 111.15 134.14 112.86 ;
   RECT 0.0 112.86 134.14 114.57 ;
   RECT 0.0 114.57 134.14 116.28 ;
   RECT 0.0 116.28 134.14 117.99 ;
   RECT 0.0 117.99 134.14 119.7 ;
   RECT 0.0 119.7 134.14 121.41 ;
   RECT 0.0 121.41 134.14 123.12 ;
   RECT 0.0 123.12 134.14 124.83 ;
   RECT 0.0 124.83 134.14 126.54 ;
   RECT 0.0 126.54 134.14 128.25 ;
   RECT 0.0 128.25 134.14 129.96 ;
   RECT 0.0 129.96 134.14 131.67 ;
   RECT 0.0 131.67 134.14 133.38 ;
   RECT 0.0 133.38 134.14 135.09 ;
   RECT 0.0 135.09 134.14 136.8 ;
   RECT 0.0 136.8 134.14 138.51 ;
   RECT 0.0 138.51 134.14 140.22 ;
   RECT 0.0 140.22 134.14 141.93 ;
   RECT 0.0 141.93 134.14 143.64 ;
   RECT 0.0 143.64 134.14 145.35 ;
   RECT 0.0 145.35 134.14 147.06 ;
   RECT 0.0 147.06 134.14 148.77 ;
   RECT 0.0 148.77 157.32 150.48 ;
   RECT 0.0 150.48 157.32 152.19 ;
   RECT 0.0 152.19 157.32 153.9 ;
   RECT 0.0 153.9 157.32 155.61 ;
   RECT 0.0 155.61 157.32 157.32 ;
   RECT 0.0 157.32 157.32 159.03 ;
   RECT 0.0 159.03 157.32 160.74 ;
   RECT 0.0 160.74 157.32 162.45 ;
   RECT 0.0 162.45 157.32 164.16 ;
   RECT 0.0 164.16 157.32 165.87 ;
   RECT 0.0 165.87 157.32 167.58 ;
   RECT 0.0 167.58 157.32 169.29 ;
   RECT 0.0 169.29 157.32 171.0 ;
   RECT 0.0 171.0 157.32 172.71 ;
   RECT 0.0 172.71 157.32 174.42 ;
   RECT 0.0 174.42 157.32 176.13 ;
   RECT 0.0 176.13 157.32 177.84 ;
   RECT 0.0 177.84 134.14 179.55 ;
   RECT 0.0 179.55 134.14 181.26 ;
   RECT 0.0 181.26 134.14 182.97 ;
   RECT 0.0 182.97 134.14 184.68 ;
   RECT 0.0 184.68 134.14 186.39 ;
   RECT 0.0 186.39 134.14 188.1 ;
   RECT 0.0 188.1 134.14 189.81 ;
   RECT 0.0 189.81 134.14 191.52 ;
   RECT 0.0 191.52 134.14 193.23 ;
   RECT 0.0 193.23 134.14 194.94 ;
   RECT 0.0 194.94 134.14 196.65 ;
   RECT 0.0 196.65 134.14 198.36 ;
   RECT 0.0 198.36 134.14 200.07 ;
   RECT 0.0 200.07 134.14 201.78 ;
   RECT 0.0 201.78 134.14 203.49 ;
   RECT 0.0 203.49 134.14 205.2 ;
   RECT 0.0 205.2 134.14 206.91 ;
   RECT 0.0 206.91 134.14 208.62 ;
   RECT 0.0 208.62 134.14 210.33 ;
   RECT 0.0 210.33 134.14 212.04 ;
   RECT 0.0 212.04 134.14 213.75 ;
   RECT 0.0 213.75 134.14 215.46 ;
   RECT 0.0 215.46 134.14 217.17 ;
   RECT 0.0 217.17 134.14 218.88 ;
   RECT 0.0 218.88 134.14 220.59 ;
   RECT 0.0 220.59 134.14 222.3 ;
   RECT 0.0 222.3 134.14 224.01 ;
   RECT 0.0 224.01 134.14 225.72 ;
   RECT 0.0 225.72 134.14 227.43 ;
   RECT 0.0 227.43 134.14 229.14 ;
   RECT 0.0 229.14 134.14 230.85 ;
   RECT 0.0 230.85 134.14 232.56 ;
   RECT 0.0 232.56 134.14 234.27 ;
   RECT 0.0 234.27 134.14 235.98 ;
   RECT 0.0 235.98 134.14 237.69 ;
   RECT 0.0 237.69 134.14 239.4 ;
   RECT 0.0 239.4 134.14 241.11 ;
   RECT 0.0 241.11 134.14 242.82 ;
   RECT 0.0 242.82 134.14 244.53 ;
   RECT 0.0 244.53 134.14 246.24 ;
   RECT 0.0 246.24 134.14 247.95 ;
   RECT 0.0 247.95 134.14 249.66 ;
   RECT 0.0 249.66 134.14 251.37 ;
   RECT 0.0 251.37 134.14 253.08 ;
   RECT 0.0 253.08 134.14 254.79 ;
   RECT 0.0 254.79 134.14 256.5 ;
   RECT 0.0 256.5 134.14 258.21 ;
   RECT 0.0 258.21 134.14 259.92 ;
   RECT 0.0 259.92 134.14 261.63 ;
   RECT 0.0 261.63 134.14 263.34 ;
   RECT 0.0 263.34 134.14 265.05 ;
   RECT 0.0 265.05 134.14 266.76 ;
   RECT 0.0 266.76 134.14 268.47 ;
   RECT 0.0 268.47 134.14 270.18 ;
   RECT 0.0 270.18 134.14 271.89 ;
   RECT 0.0 271.89 134.14 273.6 ;
   RECT 0.0 273.6 134.14 275.31 ;
   RECT 0.0 275.31 134.14 277.02 ;
   RECT 0.0 277.02 134.14 278.73 ;
   RECT 0.0 278.73 134.14 280.44 ;
   RECT 0.0 280.44 134.14 282.15 ;
   RECT 0.0 282.15 134.14 283.86 ;
   RECT 0.0 283.86 134.14 285.57 ;
   RECT 0.0 285.57 134.14 287.28 ;
   RECT 0.0 287.28 134.14 288.99 ;
   RECT 0.0 288.99 134.14 290.7 ;
   RECT 0.0 290.7 134.14 292.41 ;
   RECT 0.0 292.41 134.14 294.12 ;
   RECT 0.0 294.12 134.14 295.83 ;
   RECT 0.0 295.83 134.14 297.54 ;
   RECT 0.0 297.54 134.14 299.25 ;
   RECT 0.0 299.25 134.14 300.96 ;
   RECT 0.0 300.96 134.14 302.67 ;
   RECT 0.0 302.67 134.14 304.38 ;
   RECT 0.0 304.38 134.14 306.09 ;
   RECT 0.0 306.09 134.14 307.8 ;
   RECT 0.0 307.8 134.14 309.51 ;
   RECT 0.0 309.51 134.14 311.22 ;
   RECT 0.0 311.22 134.14 312.93 ;
   RECT 0.0 312.93 134.14 314.64 ;
   RECT 0.0 314.64 134.14 316.35 ;
   RECT 0.0 316.35 134.14 318.06 ;
   RECT 0.0 318.06 134.14 319.77 ;
   RECT 0.0 319.77 134.14 321.48 ;
   RECT 0.0 321.48 134.14 323.19 ;
   RECT 0.0 323.19 134.14 324.9 ;
   RECT 0.0 324.9 134.14 326.61 ;
   RECT 0.0 326.61 134.14 328.32 ;
   RECT 0.0 328.32 134.14 330.03 ;
   RECT 0.0 330.03 134.14 331.74 ;
  LAYER metal2 ;
   RECT 0.0 0.0 134.14 1.71 ;
   RECT 0.0 1.71 134.14 3.42 ;
   RECT 0.0 3.42 134.14 5.13 ;
   RECT 0.0 5.13 134.14 6.84 ;
   RECT 0.0 6.84 134.14 8.55 ;
   RECT 0.0 8.55 134.14 10.26 ;
   RECT 0.0 10.26 134.14 11.97 ;
   RECT 0.0 11.97 134.14 13.68 ;
   RECT 0.0 13.68 134.14 15.39 ;
   RECT 0.0 15.39 134.14 17.1 ;
   RECT 0.0 17.1 134.14 18.81 ;
   RECT 0.0 18.81 134.14 20.52 ;
   RECT 0.0 20.52 134.14 22.23 ;
   RECT 0.0 22.23 134.14 23.94 ;
   RECT 0.0 23.94 134.14 25.65 ;
   RECT 0.0 25.65 134.14 27.36 ;
   RECT 0.0 27.36 134.14 29.07 ;
   RECT 0.0 29.07 134.14 30.78 ;
   RECT 0.0 30.78 134.14 32.49 ;
   RECT 0.0 32.49 134.14 34.2 ;
   RECT 0.0 34.2 134.14 35.91 ;
   RECT 0.0 35.91 134.14 37.62 ;
   RECT 0.0 37.62 134.14 39.33 ;
   RECT 0.0 39.33 134.14 41.04 ;
   RECT 0.0 41.04 134.14 42.75 ;
   RECT 0.0 42.75 134.14 44.46 ;
   RECT 0.0 44.46 134.14 46.17 ;
   RECT 0.0 46.17 134.14 47.88 ;
   RECT 0.0 47.88 134.14 49.59 ;
   RECT 0.0 49.59 134.14 51.3 ;
   RECT 0.0 51.3 134.14 53.01 ;
   RECT 0.0 53.01 134.14 54.72 ;
   RECT 0.0 54.72 134.14 56.43 ;
   RECT 0.0 56.43 134.14 58.14 ;
   RECT 0.0 58.14 134.14 59.85 ;
   RECT 0.0 59.85 134.14 61.56 ;
   RECT 0.0 61.56 134.14 63.27 ;
   RECT 0.0 63.27 134.14 64.98 ;
   RECT 0.0 64.98 134.14 66.69 ;
   RECT 0.0 66.69 134.14 68.4 ;
   RECT 0.0 68.4 134.14 70.11 ;
   RECT 0.0 70.11 134.14 71.82 ;
   RECT 0.0 71.82 134.14 73.53 ;
   RECT 0.0 73.53 134.14 75.24 ;
   RECT 0.0 75.24 134.14 76.95 ;
   RECT 0.0 76.95 134.14 78.66 ;
   RECT 0.0 78.66 134.14 80.37 ;
   RECT 0.0 80.37 134.14 82.08 ;
   RECT 0.0 82.08 134.14 83.79 ;
   RECT 0.0 83.79 134.14 85.5 ;
   RECT 0.0 85.5 134.14 87.21 ;
   RECT 0.0 87.21 134.14 88.92 ;
   RECT 0.0 88.92 134.14 90.63 ;
   RECT 0.0 90.63 134.14 92.34 ;
   RECT 0.0 92.34 134.14 94.05 ;
   RECT 0.0 94.05 134.14 95.76 ;
   RECT 0.0 95.76 134.14 97.47 ;
   RECT 0.0 97.47 134.14 99.18 ;
   RECT 0.0 99.18 134.14 100.89 ;
   RECT 0.0 100.89 134.14 102.6 ;
   RECT 0.0 102.6 134.14 104.31 ;
   RECT 0.0 104.31 134.14 106.02 ;
   RECT 0.0 106.02 134.14 107.73 ;
   RECT 0.0 107.73 134.14 109.44 ;
   RECT 0.0 109.44 134.14 111.15 ;
   RECT 0.0 111.15 134.14 112.86 ;
   RECT 0.0 112.86 134.14 114.57 ;
   RECT 0.0 114.57 134.14 116.28 ;
   RECT 0.0 116.28 134.14 117.99 ;
   RECT 0.0 117.99 134.14 119.7 ;
   RECT 0.0 119.7 134.14 121.41 ;
   RECT 0.0 121.41 134.14 123.12 ;
   RECT 0.0 123.12 134.14 124.83 ;
   RECT 0.0 124.83 134.14 126.54 ;
   RECT 0.0 126.54 134.14 128.25 ;
   RECT 0.0 128.25 134.14 129.96 ;
   RECT 0.0 129.96 134.14 131.67 ;
   RECT 0.0 131.67 134.14 133.38 ;
   RECT 0.0 133.38 134.14 135.09 ;
   RECT 0.0 135.09 134.14 136.8 ;
   RECT 0.0 136.8 134.14 138.51 ;
   RECT 0.0 138.51 134.14 140.22 ;
   RECT 0.0 140.22 134.14 141.93 ;
   RECT 0.0 141.93 134.14 143.64 ;
   RECT 0.0 143.64 134.14 145.35 ;
   RECT 0.0 145.35 134.14 147.06 ;
   RECT 0.0 147.06 134.14 148.77 ;
   RECT 0.0 148.77 157.32 150.48 ;
   RECT 0.0 150.48 157.32 152.19 ;
   RECT 0.0 152.19 157.32 153.9 ;
   RECT 0.0 153.9 157.32 155.61 ;
   RECT 0.0 155.61 157.32 157.32 ;
   RECT 0.0 157.32 157.32 159.03 ;
   RECT 0.0 159.03 157.32 160.74 ;
   RECT 0.0 160.74 157.32 162.45 ;
   RECT 0.0 162.45 157.32 164.16 ;
   RECT 0.0 164.16 157.32 165.87 ;
   RECT 0.0 165.87 157.32 167.58 ;
   RECT 0.0 167.58 157.32 169.29 ;
   RECT 0.0 169.29 157.32 171.0 ;
   RECT 0.0 171.0 157.32 172.71 ;
   RECT 0.0 172.71 157.32 174.42 ;
   RECT 0.0 174.42 157.32 176.13 ;
   RECT 0.0 176.13 157.32 177.84 ;
   RECT 0.0 177.84 134.14 179.55 ;
   RECT 0.0 179.55 134.14 181.26 ;
   RECT 0.0 181.26 134.14 182.97 ;
   RECT 0.0 182.97 134.14 184.68 ;
   RECT 0.0 184.68 134.14 186.39 ;
   RECT 0.0 186.39 134.14 188.1 ;
   RECT 0.0 188.1 134.14 189.81 ;
   RECT 0.0 189.81 134.14 191.52 ;
   RECT 0.0 191.52 134.14 193.23 ;
   RECT 0.0 193.23 134.14 194.94 ;
   RECT 0.0 194.94 134.14 196.65 ;
   RECT 0.0 196.65 134.14 198.36 ;
   RECT 0.0 198.36 134.14 200.07 ;
   RECT 0.0 200.07 134.14 201.78 ;
   RECT 0.0 201.78 134.14 203.49 ;
   RECT 0.0 203.49 134.14 205.2 ;
   RECT 0.0 205.2 134.14 206.91 ;
   RECT 0.0 206.91 134.14 208.62 ;
   RECT 0.0 208.62 134.14 210.33 ;
   RECT 0.0 210.33 134.14 212.04 ;
   RECT 0.0 212.04 134.14 213.75 ;
   RECT 0.0 213.75 134.14 215.46 ;
   RECT 0.0 215.46 134.14 217.17 ;
   RECT 0.0 217.17 134.14 218.88 ;
   RECT 0.0 218.88 134.14 220.59 ;
   RECT 0.0 220.59 134.14 222.3 ;
   RECT 0.0 222.3 134.14 224.01 ;
   RECT 0.0 224.01 134.14 225.72 ;
   RECT 0.0 225.72 134.14 227.43 ;
   RECT 0.0 227.43 134.14 229.14 ;
   RECT 0.0 229.14 134.14 230.85 ;
   RECT 0.0 230.85 134.14 232.56 ;
   RECT 0.0 232.56 134.14 234.27 ;
   RECT 0.0 234.27 134.14 235.98 ;
   RECT 0.0 235.98 134.14 237.69 ;
   RECT 0.0 237.69 134.14 239.4 ;
   RECT 0.0 239.4 134.14 241.11 ;
   RECT 0.0 241.11 134.14 242.82 ;
   RECT 0.0 242.82 134.14 244.53 ;
   RECT 0.0 244.53 134.14 246.24 ;
   RECT 0.0 246.24 134.14 247.95 ;
   RECT 0.0 247.95 134.14 249.66 ;
   RECT 0.0 249.66 134.14 251.37 ;
   RECT 0.0 251.37 134.14 253.08 ;
   RECT 0.0 253.08 134.14 254.79 ;
   RECT 0.0 254.79 134.14 256.5 ;
   RECT 0.0 256.5 134.14 258.21 ;
   RECT 0.0 258.21 134.14 259.92 ;
   RECT 0.0 259.92 134.14 261.63 ;
   RECT 0.0 261.63 134.14 263.34 ;
   RECT 0.0 263.34 134.14 265.05 ;
   RECT 0.0 265.05 134.14 266.76 ;
   RECT 0.0 266.76 134.14 268.47 ;
   RECT 0.0 268.47 134.14 270.18 ;
   RECT 0.0 270.18 134.14 271.89 ;
   RECT 0.0 271.89 134.14 273.6 ;
   RECT 0.0 273.6 134.14 275.31 ;
   RECT 0.0 275.31 134.14 277.02 ;
   RECT 0.0 277.02 134.14 278.73 ;
   RECT 0.0 278.73 134.14 280.44 ;
   RECT 0.0 280.44 134.14 282.15 ;
   RECT 0.0 282.15 134.14 283.86 ;
   RECT 0.0 283.86 134.14 285.57 ;
   RECT 0.0 285.57 134.14 287.28 ;
   RECT 0.0 287.28 134.14 288.99 ;
   RECT 0.0 288.99 134.14 290.7 ;
   RECT 0.0 290.7 134.14 292.41 ;
   RECT 0.0 292.41 134.14 294.12 ;
   RECT 0.0 294.12 134.14 295.83 ;
   RECT 0.0 295.83 134.14 297.54 ;
   RECT 0.0 297.54 134.14 299.25 ;
   RECT 0.0 299.25 134.14 300.96 ;
   RECT 0.0 300.96 134.14 302.67 ;
   RECT 0.0 302.67 134.14 304.38 ;
   RECT 0.0 304.38 134.14 306.09 ;
   RECT 0.0 306.09 134.14 307.8 ;
   RECT 0.0 307.8 134.14 309.51 ;
   RECT 0.0 309.51 134.14 311.22 ;
   RECT 0.0 311.22 134.14 312.93 ;
   RECT 0.0 312.93 134.14 314.64 ;
   RECT 0.0 314.64 134.14 316.35 ;
   RECT 0.0 316.35 134.14 318.06 ;
   RECT 0.0 318.06 134.14 319.77 ;
   RECT 0.0 319.77 134.14 321.48 ;
   RECT 0.0 321.48 134.14 323.19 ;
   RECT 0.0 323.19 134.14 324.9 ;
   RECT 0.0 324.9 134.14 326.61 ;
   RECT 0.0 326.61 134.14 328.32 ;
   RECT 0.0 328.32 134.14 330.03 ;
   RECT 0.0 330.03 134.14 331.74 ;
  LAYER via2 ;
   RECT 0.0 0.0 134.14 1.71 ;
   RECT 0.0 1.71 134.14 3.42 ;
   RECT 0.0 3.42 134.14 5.13 ;
   RECT 0.0 5.13 134.14 6.84 ;
   RECT 0.0 6.84 134.14 8.55 ;
   RECT 0.0 8.55 134.14 10.26 ;
   RECT 0.0 10.26 134.14 11.97 ;
   RECT 0.0 11.97 134.14 13.68 ;
   RECT 0.0 13.68 134.14 15.39 ;
   RECT 0.0 15.39 134.14 17.1 ;
   RECT 0.0 17.1 134.14 18.81 ;
   RECT 0.0 18.81 134.14 20.52 ;
   RECT 0.0 20.52 134.14 22.23 ;
   RECT 0.0 22.23 134.14 23.94 ;
   RECT 0.0 23.94 134.14 25.65 ;
   RECT 0.0 25.65 134.14 27.36 ;
   RECT 0.0 27.36 134.14 29.07 ;
   RECT 0.0 29.07 134.14 30.78 ;
   RECT 0.0 30.78 134.14 32.49 ;
   RECT 0.0 32.49 134.14 34.2 ;
   RECT 0.0 34.2 134.14 35.91 ;
   RECT 0.0 35.91 134.14 37.62 ;
   RECT 0.0 37.62 134.14 39.33 ;
   RECT 0.0 39.33 134.14 41.04 ;
   RECT 0.0 41.04 134.14 42.75 ;
   RECT 0.0 42.75 134.14 44.46 ;
   RECT 0.0 44.46 134.14 46.17 ;
   RECT 0.0 46.17 134.14 47.88 ;
   RECT 0.0 47.88 134.14 49.59 ;
   RECT 0.0 49.59 134.14 51.3 ;
   RECT 0.0 51.3 134.14 53.01 ;
   RECT 0.0 53.01 134.14 54.72 ;
   RECT 0.0 54.72 134.14 56.43 ;
   RECT 0.0 56.43 134.14 58.14 ;
   RECT 0.0 58.14 134.14 59.85 ;
   RECT 0.0 59.85 134.14 61.56 ;
   RECT 0.0 61.56 134.14 63.27 ;
   RECT 0.0 63.27 134.14 64.98 ;
   RECT 0.0 64.98 134.14 66.69 ;
   RECT 0.0 66.69 134.14 68.4 ;
   RECT 0.0 68.4 134.14 70.11 ;
   RECT 0.0 70.11 134.14 71.82 ;
   RECT 0.0 71.82 134.14 73.53 ;
   RECT 0.0 73.53 134.14 75.24 ;
   RECT 0.0 75.24 134.14 76.95 ;
   RECT 0.0 76.95 134.14 78.66 ;
   RECT 0.0 78.66 134.14 80.37 ;
   RECT 0.0 80.37 134.14 82.08 ;
   RECT 0.0 82.08 134.14 83.79 ;
   RECT 0.0 83.79 134.14 85.5 ;
   RECT 0.0 85.5 134.14 87.21 ;
   RECT 0.0 87.21 134.14 88.92 ;
   RECT 0.0 88.92 134.14 90.63 ;
   RECT 0.0 90.63 134.14 92.34 ;
   RECT 0.0 92.34 134.14 94.05 ;
   RECT 0.0 94.05 134.14 95.76 ;
   RECT 0.0 95.76 134.14 97.47 ;
   RECT 0.0 97.47 134.14 99.18 ;
   RECT 0.0 99.18 134.14 100.89 ;
   RECT 0.0 100.89 134.14 102.6 ;
   RECT 0.0 102.6 134.14 104.31 ;
   RECT 0.0 104.31 134.14 106.02 ;
   RECT 0.0 106.02 134.14 107.73 ;
   RECT 0.0 107.73 134.14 109.44 ;
   RECT 0.0 109.44 134.14 111.15 ;
   RECT 0.0 111.15 134.14 112.86 ;
   RECT 0.0 112.86 134.14 114.57 ;
   RECT 0.0 114.57 134.14 116.28 ;
   RECT 0.0 116.28 134.14 117.99 ;
   RECT 0.0 117.99 134.14 119.7 ;
   RECT 0.0 119.7 134.14 121.41 ;
   RECT 0.0 121.41 134.14 123.12 ;
   RECT 0.0 123.12 134.14 124.83 ;
   RECT 0.0 124.83 134.14 126.54 ;
   RECT 0.0 126.54 134.14 128.25 ;
   RECT 0.0 128.25 134.14 129.96 ;
   RECT 0.0 129.96 134.14 131.67 ;
   RECT 0.0 131.67 134.14 133.38 ;
   RECT 0.0 133.38 134.14 135.09 ;
   RECT 0.0 135.09 134.14 136.8 ;
   RECT 0.0 136.8 134.14 138.51 ;
   RECT 0.0 138.51 134.14 140.22 ;
   RECT 0.0 140.22 134.14 141.93 ;
   RECT 0.0 141.93 134.14 143.64 ;
   RECT 0.0 143.64 134.14 145.35 ;
   RECT 0.0 145.35 134.14 147.06 ;
   RECT 0.0 147.06 134.14 148.77 ;
   RECT 0.0 148.77 157.32 150.48 ;
   RECT 0.0 150.48 157.32 152.19 ;
   RECT 0.0 152.19 157.32 153.9 ;
   RECT 0.0 153.9 157.32 155.61 ;
   RECT 0.0 155.61 157.32 157.32 ;
   RECT 0.0 157.32 157.32 159.03 ;
   RECT 0.0 159.03 157.32 160.74 ;
   RECT 0.0 160.74 157.32 162.45 ;
   RECT 0.0 162.45 157.32 164.16 ;
   RECT 0.0 164.16 157.32 165.87 ;
   RECT 0.0 165.87 157.32 167.58 ;
   RECT 0.0 167.58 157.32 169.29 ;
   RECT 0.0 169.29 157.32 171.0 ;
   RECT 0.0 171.0 157.32 172.71 ;
   RECT 0.0 172.71 157.32 174.42 ;
   RECT 0.0 174.42 157.32 176.13 ;
   RECT 0.0 176.13 157.32 177.84 ;
   RECT 0.0 177.84 134.14 179.55 ;
   RECT 0.0 179.55 134.14 181.26 ;
   RECT 0.0 181.26 134.14 182.97 ;
   RECT 0.0 182.97 134.14 184.68 ;
   RECT 0.0 184.68 134.14 186.39 ;
   RECT 0.0 186.39 134.14 188.1 ;
   RECT 0.0 188.1 134.14 189.81 ;
   RECT 0.0 189.81 134.14 191.52 ;
   RECT 0.0 191.52 134.14 193.23 ;
   RECT 0.0 193.23 134.14 194.94 ;
   RECT 0.0 194.94 134.14 196.65 ;
   RECT 0.0 196.65 134.14 198.36 ;
   RECT 0.0 198.36 134.14 200.07 ;
   RECT 0.0 200.07 134.14 201.78 ;
   RECT 0.0 201.78 134.14 203.49 ;
   RECT 0.0 203.49 134.14 205.2 ;
   RECT 0.0 205.2 134.14 206.91 ;
   RECT 0.0 206.91 134.14 208.62 ;
   RECT 0.0 208.62 134.14 210.33 ;
   RECT 0.0 210.33 134.14 212.04 ;
   RECT 0.0 212.04 134.14 213.75 ;
   RECT 0.0 213.75 134.14 215.46 ;
   RECT 0.0 215.46 134.14 217.17 ;
   RECT 0.0 217.17 134.14 218.88 ;
   RECT 0.0 218.88 134.14 220.59 ;
   RECT 0.0 220.59 134.14 222.3 ;
   RECT 0.0 222.3 134.14 224.01 ;
   RECT 0.0 224.01 134.14 225.72 ;
   RECT 0.0 225.72 134.14 227.43 ;
   RECT 0.0 227.43 134.14 229.14 ;
   RECT 0.0 229.14 134.14 230.85 ;
   RECT 0.0 230.85 134.14 232.56 ;
   RECT 0.0 232.56 134.14 234.27 ;
   RECT 0.0 234.27 134.14 235.98 ;
   RECT 0.0 235.98 134.14 237.69 ;
   RECT 0.0 237.69 134.14 239.4 ;
   RECT 0.0 239.4 134.14 241.11 ;
   RECT 0.0 241.11 134.14 242.82 ;
   RECT 0.0 242.82 134.14 244.53 ;
   RECT 0.0 244.53 134.14 246.24 ;
   RECT 0.0 246.24 134.14 247.95 ;
   RECT 0.0 247.95 134.14 249.66 ;
   RECT 0.0 249.66 134.14 251.37 ;
   RECT 0.0 251.37 134.14 253.08 ;
   RECT 0.0 253.08 134.14 254.79 ;
   RECT 0.0 254.79 134.14 256.5 ;
   RECT 0.0 256.5 134.14 258.21 ;
   RECT 0.0 258.21 134.14 259.92 ;
   RECT 0.0 259.92 134.14 261.63 ;
   RECT 0.0 261.63 134.14 263.34 ;
   RECT 0.0 263.34 134.14 265.05 ;
   RECT 0.0 265.05 134.14 266.76 ;
   RECT 0.0 266.76 134.14 268.47 ;
   RECT 0.0 268.47 134.14 270.18 ;
   RECT 0.0 270.18 134.14 271.89 ;
   RECT 0.0 271.89 134.14 273.6 ;
   RECT 0.0 273.6 134.14 275.31 ;
   RECT 0.0 275.31 134.14 277.02 ;
   RECT 0.0 277.02 134.14 278.73 ;
   RECT 0.0 278.73 134.14 280.44 ;
   RECT 0.0 280.44 134.14 282.15 ;
   RECT 0.0 282.15 134.14 283.86 ;
   RECT 0.0 283.86 134.14 285.57 ;
   RECT 0.0 285.57 134.14 287.28 ;
   RECT 0.0 287.28 134.14 288.99 ;
   RECT 0.0 288.99 134.14 290.7 ;
   RECT 0.0 290.7 134.14 292.41 ;
   RECT 0.0 292.41 134.14 294.12 ;
   RECT 0.0 294.12 134.14 295.83 ;
   RECT 0.0 295.83 134.14 297.54 ;
   RECT 0.0 297.54 134.14 299.25 ;
   RECT 0.0 299.25 134.14 300.96 ;
   RECT 0.0 300.96 134.14 302.67 ;
   RECT 0.0 302.67 134.14 304.38 ;
   RECT 0.0 304.38 134.14 306.09 ;
   RECT 0.0 306.09 134.14 307.8 ;
   RECT 0.0 307.8 134.14 309.51 ;
   RECT 0.0 309.51 134.14 311.22 ;
   RECT 0.0 311.22 134.14 312.93 ;
   RECT 0.0 312.93 134.14 314.64 ;
   RECT 0.0 314.64 134.14 316.35 ;
   RECT 0.0 316.35 134.14 318.06 ;
   RECT 0.0 318.06 134.14 319.77 ;
   RECT 0.0 319.77 134.14 321.48 ;
   RECT 0.0 321.48 134.14 323.19 ;
   RECT 0.0 323.19 134.14 324.9 ;
   RECT 0.0 324.9 134.14 326.61 ;
   RECT 0.0 326.61 134.14 328.32 ;
   RECT 0.0 328.32 134.14 330.03 ;
   RECT 0.0 330.03 134.14 331.74 ;
  LAYER metal3 ;
   RECT 0.0 0.0 134.14 1.71 ;
   RECT 0.0 1.71 134.14 3.42 ;
   RECT 0.0 3.42 134.14 5.13 ;
   RECT 0.0 5.13 134.14 6.84 ;
   RECT 0.0 6.84 134.14 8.55 ;
   RECT 0.0 8.55 134.14 10.26 ;
   RECT 0.0 10.26 134.14 11.97 ;
   RECT 0.0 11.97 134.14 13.68 ;
   RECT 0.0 13.68 134.14 15.39 ;
   RECT 0.0 15.39 134.14 17.1 ;
   RECT 0.0 17.1 134.14 18.81 ;
   RECT 0.0 18.81 134.14 20.52 ;
   RECT 0.0 20.52 134.14 22.23 ;
   RECT 0.0 22.23 134.14 23.94 ;
   RECT 0.0 23.94 134.14 25.65 ;
   RECT 0.0 25.65 134.14 27.36 ;
   RECT 0.0 27.36 134.14 29.07 ;
   RECT 0.0 29.07 134.14 30.78 ;
   RECT 0.0 30.78 134.14 32.49 ;
   RECT 0.0 32.49 134.14 34.2 ;
   RECT 0.0 34.2 134.14 35.91 ;
   RECT 0.0 35.91 134.14 37.62 ;
   RECT 0.0 37.62 134.14 39.33 ;
   RECT 0.0 39.33 134.14 41.04 ;
   RECT 0.0 41.04 134.14 42.75 ;
   RECT 0.0 42.75 134.14 44.46 ;
   RECT 0.0 44.46 134.14 46.17 ;
   RECT 0.0 46.17 134.14 47.88 ;
   RECT 0.0 47.88 134.14 49.59 ;
   RECT 0.0 49.59 134.14 51.3 ;
   RECT 0.0 51.3 134.14 53.01 ;
   RECT 0.0 53.01 134.14 54.72 ;
   RECT 0.0 54.72 134.14 56.43 ;
   RECT 0.0 56.43 134.14 58.14 ;
   RECT 0.0 58.14 134.14 59.85 ;
   RECT 0.0 59.85 134.14 61.56 ;
   RECT 0.0 61.56 134.14 63.27 ;
   RECT 0.0 63.27 134.14 64.98 ;
   RECT 0.0 64.98 134.14 66.69 ;
   RECT 0.0 66.69 134.14 68.4 ;
   RECT 0.0 68.4 134.14 70.11 ;
   RECT 0.0 70.11 134.14 71.82 ;
   RECT 0.0 71.82 134.14 73.53 ;
   RECT 0.0 73.53 134.14 75.24 ;
   RECT 0.0 75.24 134.14 76.95 ;
   RECT 0.0 76.95 134.14 78.66 ;
   RECT 0.0 78.66 134.14 80.37 ;
   RECT 0.0 80.37 134.14 82.08 ;
   RECT 0.0 82.08 134.14 83.79 ;
   RECT 0.0 83.79 134.14 85.5 ;
   RECT 0.0 85.5 134.14 87.21 ;
   RECT 0.0 87.21 134.14 88.92 ;
   RECT 0.0 88.92 134.14 90.63 ;
   RECT 0.0 90.63 134.14 92.34 ;
   RECT 0.0 92.34 134.14 94.05 ;
   RECT 0.0 94.05 134.14 95.76 ;
   RECT 0.0 95.76 134.14 97.47 ;
   RECT 0.0 97.47 134.14 99.18 ;
   RECT 0.0 99.18 134.14 100.89 ;
   RECT 0.0 100.89 134.14 102.6 ;
   RECT 0.0 102.6 134.14 104.31 ;
   RECT 0.0 104.31 134.14 106.02 ;
   RECT 0.0 106.02 134.14 107.73 ;
   RECT 0.0 107.73 134.14 109.44 ;
   RECT 0.0 109.44 134.14 111.15 ;
   RECT 0.0 111.15 134.14 112.86 ;
   RECT 0.0 112.86 134.14 114.57 ;
   RECT 0.0 114.57 134.14 116.28 ;
   RECT 0.0 116.28 134.14 117.99 ;
   RECT 0.0 117.99 134.14 119.7 ;
   RECT 0.0 119.7 134.14 121.41 ;
   RECT 0.0 121.41 134.14 123.12 ;
   RECT 0.0 123.12 134.14 124.83 ;
   RECT 0.0 124.83 134.14 126.54 ;
   RECT 0.0 126.54 134.14 128.25 ;
   RECT 0.0 128.25 134.14 129.96 ;
   RECT 0.0 129.96 134.14 131.67 ;
   RECT 0.0 131.67 134.14 133.38 ;
   RECT 0.0 133.38 134.14 135.09 ;
   RECT 0.0 135.09 134.14 136.8 ;
   RECT 0.0 136.8 134.14 138.51 ;
   RECT 0.0 138.51 134.14 140.22 ;
   RECT 0.0 140.22 134.14 141.93 ;
   RECT 0.0 141.93 134.14 143.64 ;
   RECT 0.0 143.64 134.14 145.35 ;
   RECT 0.0 145.35 134.14 147.06 ;
   RECT 0.0 147.06 134.14 148.77 ;
   RECT 0.0 148.77 157.32 150.48 ;
   RECT 0.0 150.48 157.32 152.19 ;
   RECT 0.0 152.19 157.32 153.9 ;
   RECT 0.0 153.9 157.32 155.61 ;
   RECT 0.0 155.61 157.32 157.32 ;
   RECT 0.0 157.32 157.32 159.03 ;
   RECT 0.0 159.03 157.32 160.74 ;
   RECT 0.0 160.74 157.32 162.45 ;
   RECT 0.0 162.45 157.32 164.16 ;
   RECT 0.0 164.16 157.32 165.87 ;
   RECT 0.0 165.87 157.32 167.58 ;
   RECT 0.0 167.58 157.32 169.29 ;
   RECT 0.0 169.29 157.32 171.0 ;
   RECT 0.0 171.0 157.32 172.71 ;
   RECT 0.0 172.71 157.32 174.42 ;
   RECT 0.0 174.42 157.32 176.13 ;
   RECT 0.0 176.13 157.32 177.84 ;
   RECT 0.0 177.84 134.14 179.55 ;
   RECT 0.0 179.55 134.14 181.26 ;
   RECT 0.0 181.26 134.14 182.97 ;
   RECT 0.0 182.97 134.14 184.68 ;
   RECT 0.0 184.68 134.14 186.39 ;
   RECT 0.0 186.39 134.14 188.1 ;
   RECT 0.0 188.1 134.14 189.81 ;
   RECT 0.0 189.81 134.14 191.52 ;
   RECT 0.0 191.52 134.14 193.23 ;
   RECT 0.0 193.23 134.14 194.94 ;
   RECT 0.0 194.94 134.14 196.65 ;
   RECT 0.0 196.65 134.14 198.36 ;
   RECT 0.0 198.36 134.14 200.07 ;
   RECT 0.0 200.07 134.14 201.78 ;
   RECT 0.0 201.78 134.14 203.49 ;
   RECT 0.0 203.49 134.14 205.2 ;
   RECT 0.0 205.2 134.14 206.91 ;
   RECT 0.0 206.91 134.14 208.62 ;
   RECT 0.0 208.62 134.14 210.33 ;
   RECT 0.0 210.33 134.14 212.04 ;
   RECT 0.0 212.04 134.14 213.75 ;
   RECT 0.0 213.75 134.14 215.46 ;
   RECT 0.0 215.46 134.14 217.17 ;
   RECT 0.0 217.17 134.14 218.88 ;
   RECT 0.0 218.88 134.14 220.59 ;
   RECT 0.0 220.59 134.14 222.3 ;
   RECT 0.0 222.3 134.14 224.01 ;
   RECT 0.0 224.01 134.14 225.72 ;
   RECT 0.0 225.72 134.14 227.43 ;
   RECT 0.0 227.43 134.14 229.14 ;
   RECT 0.0 229.14 134.14 230.85 ;
   RECT 0.0 230.85 134.14 232.56 ;
   RECT 0.0 232.56 134.14 234.27 ;
   RECT 0.0 234.27 134.14 235.98 ;
   RECT 0.0 235.98 134.14 237.69 ;
   RECT 0.0 237.69 134.14 239.4 ;
   RECT 0.0 239.4 134.14 241.11 ;
   RECT 0.0 241.11 134.14 242.82 ;
   RECT 0.0 242.82 134.14 244.53 ;
   RECT 0.0 244.53 134.14 246.24 ;
   RECT 0.0 246.24 134.14 247.95 ;
   RECT 0.0 247.95 134.14 249.66 ;
   RECT 0.0 249.66 134.14 251.37 ;
   RECT 0.0 251.37 134.14 253.08 ;
   RECT 0.0 253.08 134.14 254.79 ;
   RECT 0.0 254.79 134.14 256.5 ;
   RECT 0.0 256.5 134.14 258.21 ;
   RECT 0.0 258.21 134.14 259.92 ;
   RECT 0.0 259.92 134.14 261.63 ;
   RECT 0.0 261.63 134.14 263.34 ;
   RECT 0.0 263.34 134.14 265.05 ;
   RECT 0.0 265.05 134.14 266.76 ;
   RECT 0.0 266.76 134.14 268.47 ;
   RECT 0.0 268.47 134.14 270.18 ;
   RECT 0.0 270.18 134.14 271.89 ;
   RECT 0.0 271.89 134.14 273.6 ;
   RECT 0.0 273.6 134.14 275.31 ;
   RECT 0.0 275.31 134.14 277.02 ;
   RECT 0.0 277.02 134.14 278.73 ;
   RECT 0.0 278.73 134.14 280.44 ;
   RECT 0.0 280.44 134.14 282.15 ;
   RECT 0.0 282.15 134.14 283.86 ;
   RECT 0.0 283.86 134.14 285.57 ;
   RECT 0.0 285.57 134.14 287.28 ;
   RECT 0.0 287.28 134.14 288.99 ;
   RECT 0.0 288.99 134.14 290.7 ;
   RECT 0.0 290.7 134.14 292.41 ;
   RECT 0.0 292.41 134.14 294.12 ;
   RECT 0.0 294.12 134.14 295.83 ;
   RECT 0.0 295.83 134.14 297.54 ;
   RECT 0.0 297.54 134.14 299.25 ;
   RECT 0.0 299.25 134.14 300.96 ;
   RECT 0.0 300.96 134.14 302.67 ;
   RECT 0.0 302.67 134.14 304.38 ;
   RECT 0.0 304.38 134.14 306.09 ;
   RECT 0.0 306.09 134.14 307.8 ;
   RECT 0.0 307.8 134.14 309.51 ;
   RECT 0.0 309.51 134.14 311.22 ;
   RECT 0.0 311.22 134.14 312.93 ;
   RECT 0.0 312.93 134.14 314.64 ;
   RECT 0.0 314.64 134.14 316.35 ;
   RECT 0.0 316.35 134.14 318.06 ;
   RECT 0.0 318.06 134.14 319.77 ;
   RECT 0.0 319.77 134.14 321.48 ;
   RECT 0.0 321.48 134.14 323.19 ;
   RECT 0.0 323.19 134.14 324.9 ;
   RECT 0.0 324.9 134.14 326.61 ;
   RECT 0.0 326.61 134.14 328.32 ;
   RECT 0.0 328.32 134.14 330.03 ;
   RECT 0.0 330.03 134.14 331.74 ;
  LAYER via3 ;
   RECT 0.0 0.0 134.14 1.71 ;
   RECT 0.0 1.71 134.14 3.42 ;
   RECT 0.0 3.42 134.14 5.13 ;
   RECT 0.0 5.13 134.14 6.84 ;
   RECT 0.0 6.84 134.14 8.55 ;
   RECT 0.0 8.55 134.14 10.26 ;
   RECT 0.0 10.26 134.14 11.97 ;
   RECT 0.0 11.97 134.14 13.68 ;
   RECT 0.0 13.68 134.14 15.39 ;
   RECT 0.0 15.39 134.14 17.1 ;
   RECT 0.0 17.1 134.14 18.81 ;
   RECT 0.0 18.81 134.14 20.52 ;
   RECT 0.0 20.52 134.14 22.23 ;
   RECT 0.0 22.23 134.14 23.94 ;
   RECT 0.0 23.94 134.14 25.65 ;
   RECT 0.0 25.65 134.14 27.36 ;
   RECT 0.0 27.36 134.14 29.07 ;
   RECT 0.0 29.07 134.14 30.78 ;
   RECT 0.0 30.78 134.14 32.49 ;
   RECT 0.0 32.49 134.14 34.2 ;
   RECT 0.0 34.2 134.14 35.91 ;
   RECT 0.0 35.91 134.14 37.62 ;
   RECT 0.0 37.62 134.14 39.33 ;
   RECT 0.0 39.33 134.14 41.04 ;
   RECT 0.0 41.04 134.14 42.75 ;
   RECT 0.0 42.75 134.14 44.46 ;
   RECT 0.0 44.46 134.14 46.17 ;
   RECT 0.0 46.17 134.14 47.88 ;
   RECT 0.0 47.88 134.14 49.59 ;
   RECT 0.0 49.59 134.14 51.3 ;
   RECT 0.0 51.3 134.14 53.01 ;
   RECT 0.0 53.01 134.14 54.72 ;
   RECT 0.0 54.72 134.14 56.43 ;
   RECT 0.0 56.43 134.14 58.14 ;
   RECT 0.0 58.14 134.14 59.85 ;
   RECT 0.0 59.85 134.14 61.56 ;
   RECT 0.0 61.56 134.14 63.27 ;
   RECT 0.0 63.27 134.14 64.98 ;
   RECT 0.0 64.98 134.14 66.69 ;
   RECT 0.0 66.69 134.14 68.4 ;
   RECT 0.0 68.4 134.14 70.11 ;
   RECT 0.0 70.11 134.14 71.82 ;
   RECT 0.0 71.82 134.14 73.53 ;
   RECT 0.0 73.53 134.14 75.24 ;
   RECT 0.0 75.24 134.14 76.95 ;
   RECT 0.0 76.95 134.14 78.66 ;
   RECT 0.0 78.66 134.14 80.37 ;
   RECT 0.0 80.37 134.14 82.08 ;
   RECT 0.0 82.08 134.14 83.79 ;
   RECT 0.0 83.79 134.14 85.5 ;
   RECT 0.0 85.5 134.14 87.21 ;
   RECT 0.0 87.21 134.14 88.92 ;
   RECT 0.0 88.92 134.14 90.63 ;
   RECT 0.0 90.63 134.14 92.34 ;
   RECT 0.0 92.34 134.14 94.05 ;
   RECT 0.0 94.05 134.14 95.76 ;
   RECT 0.0 95.76 134.14 97.47 ;
   RECT 0.0 97.47 134.14 99.18 ;
   RECT 0.0 99.18 134.14 100.89 ;
   RECT 0.0 100.89 134.14 102.6 ;
   RECT 0.0 102.6 134.14 104.31 ;
   RECT 0.0 104.31 134.14 106.02 ;
   RECT 0.0 106.02 134.14 107.73 ;
   RECT 0.0 107.73 134.14 109.44 ;
   RECT 0.0 109.44 134.14 111.15 ;
   RECT 0.0 111.15 134.14 112.86 ;
   RECT 0.0 112.86 134.14 114.57 ;
   RECT 0.0 114.57 134.14 116.28 ;
   RECT 0.0 116.28 134.14 117.99 ;
   RECT 0.0 117.99 134.14 119.7 ;
   RECT 0.0 119.7 134.14 121.41 ;
   RECT 0.0 121.41 134.14 123.12 ;
   RECT 0.0 123.12 134.14 124.83 ;
   RECT 0.0 124.83 134.14 126.54 ;
   RECT 0.0 126.54 134.14 128.25 ;
   RECT 0.0 128.25 134.14 129.96 ;
   RECT 0.0 129.96 134.14 131.67 ;
   RECT 0.0 131.67 134.14 133.38 ;
   RECT 0.0 133.38 134.14 135.09 ;
   RECT 0.0 135.09 134.14 136.8 ;
   RECT 0.0 136.8 134.14 138.51 ;
   RECT 0.0 138.51 134.14 140.22 ;
   RECT 0.0 140.22 134.14 141.93 ;
   RECT 0.0 141.93 134.14 143.64 ;
   RECT 0.0 143.64 134.14 145.35 ;
   RECT 0.0 145.35 134.14 147.06 ;
   RECT 0.0 147.06 134.14 148.77 ;
   RECT 0.0 148.77 157.32 150.48 ;
   RECT 0.0 150.48 157.32 152.19 ;
   RECT 0.0 152.19 157.32 153.9 ;
   RECT 0.0 153.9 157.32 155.61 ;
   RECT 0.0 155.61 157.32 157.32 ;
   RECT 0.0 157.32 157.32 159.03 ;
   RECT 0.0 159.03 157.32 160.74 ;
   RECT 0.0 160.74 157.32 162.45 ;
   RECT 0.0 162.45 157.32 164.16 ;
   RECT 0.0 164.16 157.32 165.87 ;
   RECT 0.0 165.87 157.32 167.58 ;
   RECT 0.0 167.58 157.32 169.29 ;
   RECT 0.0 169.29 157.32 171.0 ;
   RECT 0.0 171.0 157.32 172.71 ;
   RECT 0.0 172.71 157.32 174.42 ;
   RECT 0.0 174.42 157.32 176.13 ;
   RECT 0.0 176.13 157.32 177.84 ;
   RECT 0.0 177.84 134.14 179.55 ;
   RECT 0.0 179.55 134.14 181.26 ;
   RECT 0.0 181.26 134.14 182.97 ;
   RECT 0.0 182.97 134.14 184.68 ;
   RECT 0.0 184.68 134.14 186.39 ;
   RECT 0.0 186.39 134.14 188.1 ;
   RECT 0.0 188.1 134.14 189.81 ;
   RECT 0.0 189.81 134.14 191.52 ;
   RECT 0.0 191.52 134.14 193.23 ;
   RECT 0.0 193.23 134.14 194.94 ;
   RECT 0.0 194.94 134.14 196.65 ;
   RECT 0.0 196.65 134.14 198.36 ;
   RECT 0.0 198.36 134.14 200.07 ;
   RECT 0.0 200.07 134.14 201.78 ;
   RECT 0.0 201.78 134.14 203.49 ;
   RECT 0.0 203.49 134.14 205.2 ;
   RECT 0.0 205.2 134.14 206.91 ;
   RECT 0.0 206.91 134.14 208.62 ;
   RECT 0.0 208.62 134.14 210.33 ;
   RECT 0.0 210.33 134.14 212.04 ;
   RECT 0.0 212.04 134.14 213.75 ;
   RECT 0.0 213.75 134.14 215.46 ;
   RECT 0.0 215.46 134.14 217.17 ;
   RECT 0.0 217.17 134.14 218.88 ;
   RECT 0.0 218.88 134.14 220.59 ;
   RECT 0.0 220.59 134.14 222.3 ;
   RECT 0.0 222.3 134.14 224.01 ;
   RECT 0.0 224.01 134.14 225.72 ;
   RECT 0.0 225.72 134.14 227.43 ;
   RECT 0.0 227.43 134.14 229.14 ;
   RECT 0.0 229.14 134.14 230.85 ;
   RECT 0.0 230.85 134.14 232.56 ;
   RECT 0.0 232.56 134.14 234.27 ;
   RECT 0.0 234.27 134.14 235.98 ;
   RECT 0.0 235.98 134.14 237.69 ;
   RECT 0.0 237.69 134.14 239.4 ;
   RECT 0.0 239.4 134.14 241.11 ;
   RECT 0.0 241.11 134.14 242.82 ;
   RECT 0.0 242.82 134.14 244.53 ;
   RECT 0.0 244.53 134.14 246.24 ;
   RECT 0.0 246.24 134.14 247.95 ;
   RECT 0.0 247.95 134.14 249.66 ;
   RECT 0.0 249.66 134.14 251.37 ;
   RECT 0.0 251.37 134.14 253.08 ;
   RECT 0.0 253.08 134.14 254.79 ;
   RECT 0.0 254.79 134.14 256.5 ;
   RECT 0.0 256.5 134.14 258.21 ;
   RECT 0.0 258.21 134.14 259.92 ;
   RECT 0.0 259.92 134.14 261.63 ;
   RECT 0.0 261.63 134.14 263.34 ;
   RECT 0.0 263.34 134.14 265.05 ;
   RECT 0.0 265.05 134.14 266.76 ;
   RECT 0.0 266.76 134.14 268.47 ;
   RECT 0.0 268.47 134.14 270.18 ;
   RECT 0.0 270.18 134.14 271.89 ;
   RECT 0.0 271.89 134.14 273.6 ;
   RECT 0.0 273.6 134.14 275.31 ;
   RECT 0.0 275.31 134.14 277.02 ;
   RECT 0.0 277.02 134.14 278.73 ;
   RECT 0.0 278.73 134.14 280.44 ;
   RECT 0.0 280.44 134.14 282.15 ;
   RECT 0.0 282.15 134.14 283.86 ;
   RECT 0.0 283.86 134.14 285.57 ;
   RECT 0.0 285.57 134.14 287.28 ;
   RECT 0.0 287.28 134.14 288.99 ;
   RECT 0.0 288.99 134.14 290.7 ;
   RECT 0.0 290.7 134.14 292.41 ;
   RECT 0.0 292.41 134.14 294.12 ;
   RECT 0.0 294.12 134.14 295.83 ;
   RECT 0.0 295.83 134.14 297.54 ;
   RECT 0.0 297.54 134.14 299.25 ;
   RECT 0.0 299.25 134.14 300.96 ;
   RECT 0.0 300.96 134.14 302.67 ;
   RECT 0.0 302.67 134.14 304.38 ;
   RECT 0.0 304.38 134.14 306.09 ;
   RECT 0.0 306.09 134.14 307.8 ;
   RECT 0.0 307.8 134.14 309.51 ;
   RECT 0.0 309.51 134.14 311.22 ;
   RECT 0.0 311.22 134.14 312.93 ;
   RECT 0.0 312.93 134.14 314.64 ;
   RECT 0.0 314.64 134.14 316.35 ;
   RECT 0.0 316.35 134.14 318.06 ;
   RECT 0.0 318.06 134.14 319.77 ;
   RECT 0.0 319.77 134.14 321.48 ;
   RECT 0.0 321.48 134.14 323.19 ;
   RECT 0.0 323.19 134.14 324.9 ;
   RECT 0.0 324.9 134.14 326.61 ;
   RECT 0.0 326.61 134.14 328.32 ;
   RECT 0.0 328.32 134.14 330.03 ;
   RECT 0.0 330.03 134.14 331.74 ;
  LAYER metal4 ;
   RECT 0.0 0.0 134.14 1.71 ;
   RECT 0.0 1.71 134.14 3.42 ;
   RECT 0.0 3.42 134.14 5.13 ;
   RECT 0.0 5.13 134.14 6.84 ;
   RECT 0.0 6.84 134.14 8.55 ;
   RECT 0.0 8.55 134.14 10.26 ;
   RECT 0.0 10.26 134.14 11.97 ;
   RECT 0.0 11.97 134.14 13.68 ;
   RECT 0.0 13.68 134.14 15.39 ;
   RECT 0.0 15.39 134.14 17.1 ;
   RECT 0.0 17.1 134.14 18.81 ;
   RECT 0.0 18.81 134.14 20.52 ;
   RECT 0.0 20.52 134.14 22.23 ;
   RECT 0.0 22.23 134.14 23.94 ;
   RECT 0.0 23.94 134.14 25.65 ;
   RECT 0.0 25.65 134.14 27.36 ;
   RECT 0.0 27.36 134.14 29.07 ;
   RECT 0.0 29.07 134.14 30.78 ;
   RECT 0.0 30.78 134.14 32.49 ;
   RECT 0.0 32.49 134.14 34.2 ;
   RECT 0.0 34.2 134.14 35.91 ;
   RECT 0.0 35.91 134.14 37.62 ;
   RECT 0.0 37.62 134.14 39.33 ;
   RECT 0.0 39.33 134.14 41.04 ;
   RECT 0.0 41.04 134.14 42.75 ;
   RECT 0.0 42.75 134.14 44.46 ;
   RECT 0.0 44.46 134.14 46.17 ;
   RECT 0.0 46.17 134.14 47.88 ;
   RECT 0.0 47.88 134.14 49.59 ;
   RECT 0.0 49.59 134.14 51.3 ;
   RECT 0.0 51.3 134.14 53.01 ;
   RECT 0.0 53.01 134.14 54.72 ;
   RECT 0.0 54.72 134.14 56.43 ;
   RECT 0.0 56.43 134.14 58.14 ;
   RECT 0.0 58.14 134.14 59.85 ;
   RECT 0.0 59.85 134.14 61.56 ;
   RECT 0.0 61.56 134.14 63.27 ;
   RECT 0.0 63.27 134.14 64.98 ;
   RECT 0.0 64.98 134.14 66.69 ;
   RECT 0.0 66.69 134.14 68.4 ;
   RECT 0.0 68.4 134.14 70.11 ;
   RECT 0.0 70.11 134.14 71.82 ;
   RECT 0.0 71.82 134.14 73.53 ;
   RECT 0.0 73.53 134.14 75.24 ;
   RECT 0.0 75.24 134.14 76.95 ;
   RECT 0.0 76.95 134.14 78.66 ;
   RECT 0.0 78.66 134.14 80.37 ;
   RECT 0.0 80.37 134.14 82.08 ;
   RECT 0.0 82.08 134.14 83.79 ;
   RECT 0.0 83.79 134.14 85.5 ;
   RECT 0.0 85.5 134.14 87.21 ;
   RECT 0.0 87.21 134.14 88.92 ;
   RECT 0.0 88.92 134.14 90.63 ;
   RECT 0.0 90.63 134.14 92.34 ;
   RECT 0.0 92.34 134.14 94.05 ;
   RECT 0.0 94.05 134.14 95.76 ;
   RECT 0.0 95.76 134.14 97.47 ;
   RECT 0.0 97.47 134.14 99.18 ;
   RECT 0.0 99.18 134.14 100.89 ;
   RECT 0.0 100.89 134.14 102.6 ;
   RECT 0.0 102.6 134.14 104.31 ;
   RECT 0.0 104.31 134.14 106.02 ;
   RECT 0.0 106.02 134.14 107.73 ;
   RECT 0.0 107.73 134.14 109.44 ;
   RECT 0.0 109.44 134.14 111.15 ;
   RECT 0.0 111.15 134.14 112.86 ;
   RECT 0.0 112.86 134.14 114.57 ;
   RECT 0.0 114.57 134.14 116.28 ;
   RECT 0.0 116.28 134.14 117.99 ;
   RECT 0.0 117.99 134.14 119.7 ;
   RECT 0.0 119.7 134.14 121.41 ;
   RECT 0.0 121.41 134.14 123.12 ;
   RECT 0.0 123.12 134.14 124.83 ;
   RECT 0.0 124.83 134.14 126.54 ;
   RECT 0.0 126.54 134.14 128.25 ;
   RECT 0.0 128.25 134.14 129.96 ;
   RECT 0.0 129.96 134.14 131.67 ;
   RECT 0.0 131.67 134.14 133.38 ;
   RECT 0.0 133.38 134.14 135.09 ;
   RECT 0.0 135.09 134.14 136.8 ;
   RECT 0.0 136.8 134.14 138.51 ;
   RECT 0.0 138.51 134.14 140.22 ;
   RECT 0.0 140.22 134.14 141.93 ;
   RECT 0.0 141.93 134.14 143.64 ;
   RECT 0.0 143.64 134.14 145.35 ;
   RECT 0.0 145.35 134.14 147.06 ;
   RECT 0.0 147.06 134.14 148.77 ;
   RECT 0.0 148.77 157.32 150.48 ;
   RECT 0.0 150.48 157.32 152.19 ;
   RECT 0.0 152.19 157.32 153.9 ;
   RECT 0.0 153.9 157.32 155.61 ;
   RECT 0.0 155.61 157.32 157.32 ;
   RECT 0.0 157.32 157.32 159.03 ;
   RECT 0.0 159.03 157.32 160.74 ;
   RECT 0.0 160.74 157.32 162.45 ;
   RECT 0.0 162.45 157.32 164.16 ;
   RECT 0.0 164.16 157.32 165.87 ;
   RECT 0.0 165.87 157.32 167.58 ;
   RECT 0.0 167.58 157.32 169.29 ;
   RECT 0.0 169.29 157.32 171.0 ;
   RECT 0.0 171.0 157.32 172.71 ;
   RECT 0.0 172.71 157.32 174.42 ;
   RECT 0.0 174.42 157.32 176.13 ;
   RECT 0.0 176.13 157.32 177.84 ;
   RECT 0.0 177.84 134.14 179.55 ;
   RECT 0.0 179.55 134.14 181.26 ;
   RECT 0.0 181.26 134.14 182.97 ;
   RECT 0.0 182.97 134.14 184.68 ;
   RECT 0.0 184.68 134.14 186.39 ;
   RECT 0.0 186.39 134.14 188.1 ;
   RECT 0.0 188.1 134.14 189.81 ;
   RECT 0.0 189.81 134.14 191.52 ;
   RECT 0.0 191.52 134.14 193.23 ;
   RECT 0.0 193.23 134.14 194.94 ;
   RECT 0.0 194.94 134.14 196.65 ;
   RECT 0.0 196.65 134.14 198.36 ;
   RECT 0.0 198.36 134.14 200.07 ;
   RECT 0.0 200.07 134.14 201.78 ;
   RECT 0.0 201.78 134.14 203.49 ;
   RECT 0.0 203.49 134.14 205.2 ;
   RECT 0.0 205.2 134.14 206.91 ;
   RECT 0.0 206.91 134.14 208.62 ;
   RECT 0.0 208.62 134.14 210.33 ;
   RECT 0.0 210.33 134.14 212.04 ;
   RECT 0.0 212.04 134.14 213.75 ;
   RECT 0.0 213.75 134.14 215.46 ;
   RECT 0.0 215.46 134.14 217.17 ;
   RECT 0.0 217.17 134.14 218.88 ;
   RECT 0.0 218.88 134.14 220.59 ;
   RECT 0.0 220.59 134.14 222.3 ;
   RECT 0.0 222.3 134.14 224.01 ;
   RECT 0.0 224.01 134.14 225.72 ;
   RECT 0.0 225.72 134.14 227.43 ;
   RECT 0.0 227.43 134.14 229.14 ;
   RECT 0.0 229.14 134.14 230.85 ;
   RECT 0.0 230.85 134.14 232.56 ;
   RECT 0.0 232.56 134.14 234.27 ;
   RECT 0.0 234.27 134.14 235.98 ;
   RECT 0.0 235.98 134.14 237.69 ;
   RECT 0.0 237.69 134.14 239.4 ;
   RECT 0.0 239.4 134.14 241.11 ;
   RECT 0.0 241.11 134.14 242.82 ;
   RECT 0.0 242.82 134.14 244.53 ;
   RECT 0.0 244.53 134.14 246.24 ;
   RECT 0.0 246.24 134.14 247.95 ;
   RECT 0.0 247.95 134.14 249.66 ;
   RECT 0.0 249.66 134.14 251.37 ;
   RECT 0.0 251.37 134.14 253.08 ;
   RECT 0.0 253.08 134.14 254.79 ;
   RECT 0.0 254.79 134.14 256.5 ;
   RECT 0.0 256.5 134.14 258.21 ;
   RECT 0.0 258.21 134.14 259.92 ;
   RECT 0.0 259.92 134.14 261.63 ;
   RECT 0.0 261.63 134.14 263.34 ;
   RECT 0.0 263.34 134.14 265.05 ;
   RECT 0.0 265.05 134.14 266.76 ;
   RECT 0.0 266.76 134.14 268.47 ;
   RECT 0.0 268.47 134.14 270.18 ;
   RECT 0.0 270.18 134.14 271.89 ;
   RECT 0.0 271.89 134.14 273.6 ;
   RECT 0.0 273.6 134.14 275.31 ;
   RECT 0.0 275.31 134.14 277.02 ;
   RECT 0.0 277.02 134.14 278.73 ;
   RECT 0.0 278.73 134.14 280.44 ;
   RECT 0.0 280.44 134.14 282.15 ;
   RECT 0.0 282.15 134.14 283.86 ;
   RECT 0.0 283.86 134.14 285.57 ;
   RECT 0.0 285.57 134.14 287.28 ;
   RECT 0.0 287.28 134.14 288.99 ;
   RECT 0.0 288.99 134.14 290.7 ;
   RECT 0.0 290.7 134.14 292.41 ;
   RECT 0.0 292.41 134.14 294.12 ;
   RECT 0.0 294.12 134.14 295.83 ;
   RECT 0.0 295.83 134.14 297.54 ;
   RECT 0.0 297.54 134.14 299.25 ;
   RECT 0.0 299.25 134.14 300.96 ;
   RECT 0.0 300.96 134.14 302.67 ;
   RECT 0.0 302.67 134.14 304.38 ;
   RECT 0.0 304.38 134.14 306.09 ;
   RECT 0.0 306.09 134.14 307.8 ;
   RECT 0.0 307.8 134.14 309.51 ;
   RECT 0.0 309.51 134.14 311.22 ;
   RECT 0.0 311.22 134.14 312.93 ;
   RECT 0.0 312.93 134.14 314.64 ;
   RECT 0.0 314.64 134.14 316.35 ;
   RECT 0.0 316.35 134.14 318.06 ;
   RECT 0.0 318.06 134.14 319.77 ;
   RECT 0.0 319.77 134.14 321.48 ;
   RECT 0.0 321.48 134.14 323.19 ;
   RECT 0.0 323.19 134.14 324.9 ;
   RECT 0.0 324.9 134.14 326.61 ;
   RECT 0.0 326.61 134.14 328.32 ;
   RECT 0.0 328.32 134.14 330.03 ;
   RECT 0.0 330.03 134.14 331.74 ;
 END
END block_414x1746_310

MACRO block_341x369_75
 CLASS BLOCK ;
 FOREIGN block_341x369_75 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 129.58 BY 70.11 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 20.235 126.445 20.805 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 26.695 126.445 27.265 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 6.935 3.325 7.505 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 9.215 3.325 9.785 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 10.735 3.325 11.305 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 13.015 3.325 13.585 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 13.395 4.085 13.965 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 13.775 3.325 14.345 ;
  END
 END o7
 PIN o8
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 15.295 3.325 15.865 ;
  END
 END o8
 PIN o9
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 16.055 3.325 16.625 ;
  END
 END o9
 PIN o10
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 16.815 3.325 17.385 ;
  END
 END o10
 PIN o11
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 12.635 4.085 13.205 ;
  END
 END o11
 PIN o12
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 19.855 3.325 20.425 ;
  END
 END o12
 PIN o13
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 20.615 3.325 21.185 ;
  END
 END o13
 PIN o14
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 21.375 3.325 21.945 ;
  END
 END o14
 PIN o15
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 22.135 3.325 22.705 ;
  END
 END o15
 PIN o16
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 22.895 3.325 23.465 ;
  END
 END o16
 PIN o17
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 18.335 3.325 18.905 ;
  END
 END o17
 PIN o18
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 25.935 3.325 26.505 ;
  END
 END o18
 PIN o19
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 26.695 3.325 27.265 ;
  END
 END o19
 PIN o20
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 27.455 3.325 28.025 ;
  END
 END o20
 PIN o21
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 28.975 3.325 29.545 ;
  END
 END o21
 PIN o22
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 29.735 3.325 30.305 ;
  END
 END o22
 PIN o23
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 25.175 3.325 25.745 ;
  END
 END o23
 PIN o24
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 32.015 3.325 32.585 ;
  END
 END o24
 PIN o25
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 33.535 3.325 34.105 ;
  END
 END o25
 PIN o26
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 34.295 3.325 34.865 ;
  END
 END o26
 PIN o27
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 35.055 3.325 35.625 ;
  END
 END o27
 PIN o28
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 35.815 3.325 36.385 ;
  END
 END o28
 PIN o29
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 31.255 3.325 31.825 ;
  END
 END o29
 PIN o30
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 38.095 126.445 38.665 ;
  END
 END o30
 PIN o31
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 38.855 126.445 39.425 ;
  END
 END o31
 PIN o32
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 39.615 126.445 40.185 ;
  END
 END o32
 PIN o33
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 21.755 126.445 22.325 ;
  END
 END o33
 PIN o34
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 31.255 126.445 31.825 ;
  END
 END o34
 PIN o35
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 32.015 126.445 32.585 ;
  END
 END o35
 PIN o36
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 33.535 126.445 34.105 ;
  END
 END o36
 PIN o37
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 30.495 126.445 31.065 ;
  END
 END o37
 PIN o38
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 28.975 126.445 29.545 ;
  END
 END o38
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 35.815 126.445 36.385 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 43.035 126.445 43.605 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 32.395 125.685 32.965 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 35.435 125.685 36.005 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 36.955 126.445 37.525 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 36.575 125.685 37.145 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 33.915 125.685 34.485 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 30.115 125.685 30.685 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 40.375 3.325 40.945 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 8.455 3.325 9.025 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 25.935 126.445 26.505 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 25.175 126.445 25.745 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 24.415 126.445 24.985 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 34.675 126.445 35.245 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 30.875 125.685 31.445 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 40.755 126.445 41.325 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 27.455 126.445 28.025 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 38.475 125.685 39.045 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 39.995 125.685 40.565 ;
  END
 END i18
 PIN i19
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 39.235 125.685 39.805 ;
  END
 END i19
 PIN i20
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 124.355 40.375 124.925 40.945 ;
  END
 END i20
 PIN i21
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 8.455 126.445 9.025 ;
  END
 END i21
 PIN i22
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 9.215 126.445 9.785 ;
  END
 END i22
 PIN i23
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 10.735 126.445 11.305 ;
  END
 END i23
 PIN i24
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 11.495 126.445 12.065 ;
  END
 END i24
 PIN i25
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 12.255 126.445 12.825 ;
  END
 END i25
 PIN i26
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 13.015 126.445 13.585 ;
  END
 END i26
 PIN i27
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 8.075 125.685 8.645 ;
  END
 END i27
 PIN i28
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 7.695 126.445 8.265 ;
  END
 END i28
 PIN i29
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 7.315 125.685 7.885 ;
  END
 END i29
 PIN i30
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 6.935 126.445 7.505 ;
  END
 END i30
 PIN i31
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 6.555 125.685 7.125 ;
  END
 END i31
 PIN i32
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 13.775 126.445 14.345 ;
  END
 END i32
 PIN i33
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 15.295 126.445 15.865 ;
  END
 END i33
 PIN i34
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 16.055 126.445 16.625 ;
  END
 END i34
 PIN i35
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 16.815 126.445 17.385 ;
  END
 END i35
 OBS
  LAYER metal1 ;
   RECT 0 0 129.58 70.11 ;
  LAYER via1 ;
   RECT 0 0 129.58 70.11 ;
  LAYER metal2 ;
   RECT 0 0 129.58 70.11 ;
  LAYER via2 ;
   RECT 0 0 129.58 70.11 ;
  LAYER metal3 ;
   RECT 0 0 129.58 70.11 ;
  LAYER via3 ;
   RECT 0 0 129.58 70.11 ;
  LAYER metal4 ;
   RECT 0 0 129.58 70.11 ;
 END
END block_341x369_75

MACRO block_533x1125_87
 CLASS BLOCK ;
 FOREIGN block_533x1125_87 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 202.54 BY 213.75 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 8.455 176.225 9.025 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 24.795 176.225 25.365 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 41.135 176.225 41.705 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 75.715 176.225 76.285 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 92.055 176.225 92.625 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 136.515 176.225 137.085 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 152.855 176.225 153.425 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 187.435 176.225 188.005 ;
  END
 END o7
 PIN o8
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 203.775 176.225 204.345 ;
  END
 END o8
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.835 103.075 199.405 103.645 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.835 120.175 199.405 120.745 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.835 108.395 199.405 108.965 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.835 112.765 199.405 113.335 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.835 115.615 199.405 116.185 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.075 103.455 198.645 104.025 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.075 102.695 198.645 103.265 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.835 102.315 199.405 102.885 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.835 112.005 199.405 112.575 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.835 125.115 199.405 125.685 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.075 119.795 198.645 120.365 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.835 119.415 199.405 119.985 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.835 121.505 199.405 122.075 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.835 123.975 199.405 124.545 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.075 125.495 198.645 126.065 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 188.955 101.935 189.525 102.505 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 188.955 115.235 189.525 115.805 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 6.745 176.225 7.315 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 23.085 176.225 23.655 ;
  END
 END i18
 PIN i19
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 39.425 176.225 39.995 ;
  END
 END i19
 PIN i20
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 74.005 176.225 74.575 ;
  END
 END i20
 PIN i21
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 90.345 176.225 90.915 ;
  END
 END i21
 PIN i22
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 138.225 176.225 138.795 ;
  END
 END i22
 PIN i23
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 154.565 176.225 155.135 ;
  END
 END i23
 PIN i24
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 189.145 176.225 189.715 ;
  END
 END i24
 PIN i25
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 205.485 176.225 206.055 ;
  END
 END i25
 PIN i26
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 25.365 175.465 25.935 ;
  END
 END i26
 PIN i27
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 29.355 176.225 29.925 ;
  END
 END i27
 PIN i28
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 33.535 176.225 34.105 ;
  END
 END i28
 PIN i29
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 17.195 176.225 17.765 ;
  END
 END i29
 PIN i30
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 92.625 175.465 93.195 ;
  END
 END i30
 PIN i31
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 96.615 176.225 97.185 ;
  END
 END i31
 PIN i32
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 100.795 176.225 101.365 ;
  END
 END i32
 PIN i33
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 84.455 176.225 85.025 ;
  END
 END i33
 PIN i34
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 135.945 175.465 136.515 ;
  END
 END i34
 PIN i35
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 131.955 176.225 132.525 ;
  END
 END i35
 PIN i36
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 127.775 176.225 128.345 ;
  END
 END i36
 PIN i37
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 144.115 176.225 144.685 ;
  END
 END i37
 PIN i38
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 203.205 175.465 203.775 ;
  END
 END i38
 PIN i39
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 199.215 176.225 199.785 ;
  END
 END i39
 PIN i40
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 195.035 176.225 195.605 ;
  END
 END i40
 PIN i41
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 191.045 176.225 191.615 ;
  END
 END i41
 PIN i42
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 21.185 176.225 21.755 ;
  END
 END i42
 PIN i43
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 88.445 176.225 89.015 ;
  END
 END i43
 PIN i44
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 140.125 176.225 140.695 ;
  END
 END i44
 PIN i45
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 207.385 176.225 207.955 ;
  END
 END i45
 PIN i46
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 184.015 101.935 184.585 102.505 ;
  END
 END i46
 PIN i47
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 184.015 115.235 184.585 115.805 ;
  END
 END i47
 PIN i48
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 7.315 175.465 7.885 ;
  END
 END i48
 PIN i49
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 23.655 175.465 24.225 ;
  END
 END i49
 PIN i50
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 39.995 175.465 40.565 ;
  END
 END i50
 PIN i51
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 74.575 175.465 75.145 ;
  END
 END i51
 PIN i52
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 90.915 175.465 91.485 ;
  END
 END i52
 PIN i53
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 137.655 175.465 138.225 ;
  END
 END i53
 PIN i54
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 153.995 175.465 154.565 ;
  END
 END i54
 PIN i55
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 188.575 175.465 189.145 ;
  END
 END i55
 PIN i56
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 204.915 175.465 205.485 ;
  END
 END i56
 PIN i57
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.835 109.535 199.405 110.105 ;
  END
 END i57
 PIN i58
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.075 109.915 198.645 110.485 ;
  END
 END i58
 PIN i59
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 7.885 174.705 8.455 ;
  END
 END i59
 PIN i60
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 24.225 174.705 24.795 ;
  END
 END i60
 PIN i61
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 40.565 174.705 41.135 ;
  END
 END i61
 PIN i62
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 75.145 174.705 75.715 ;
  END
 END i62
 PIN i63
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 91.485 174.705 92.055 ;
  END
 END i63
 PIN i64
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 137.085 174.705 137.655 ;
  END
 END i64
 PIN i65
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 153.425 174.705 153.995 ;
  END
 END i65
 PIN i66
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 188.005 174.705 188.575 ;
  END
 END i66
 PIN i67
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 204.345 174.705 204.915 ;
  END
 END i67
 PIN i68
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 197.695 101.935 198.265 102.505 ;
  END
 END i68
 PIN i69
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 196.555 101.935 197.125 102.505 ;
  END
 END i69
 PIN i70
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 195.035 101.935 195.605 102.505 ;
  END
 END i70
 PIN i71
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 193.135 101.935 193.705 102.505 ;
  END
 END i71
 PIN i72
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 191.995 101.935 192.565 102.505 ;
  END
 END i72
 PIN i73
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 197.695 115.235 198.265 115.805 ;
  END
 END i73
 PIN i74
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 196.555 115.235 197.125 115.805 ;
  END
 END i74
 PIN i75
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 195.035 115.235 195.605 115.805 ;
  END
 END i75
 PIN i76
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 193.135 115.235 193.705 115.805 ;
  END
 END i76
 PIN i77
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 191.995 115.235 192.565 115.805 ;
  END
 END i77
 OBS
  LAYER metal1 ;
   RECT 0.0 0.0 179.36 1.71 ;
   RECT 0.0 1.71 179.36 3.42 ;
   RECT 0.0 3.42 179.36 5.13 ;
   RECT 0.0 5.13 179.36 6.84 ;
   RECT 0.0 6.84 179.36 8.55 ;
   RECT 0.0 8.55 179.36 10.26 ;
   RECT 0.0 10.26 179.36 11.97 ;
   RECT 0.0 11.97 179.36 13.68 ;
   RECT 0.0 13.68 179.36 15.39 ;
   RECT 0.0 15.39 179.36 17.1 ;
   RECT 0.0 17.1 179.36 18.81 ;
   RECT 0.0 18.81 179.36 20.52 ;
   RECT 0.0 20.52 179.36 22.23 ;
   RECT 0.0 22.23 179.36 23.94 ;
   RECT 0.0 23.94 179.36 25.65 ;
   RECT 0.0 25.65 179.36 27.36 ;
   RECT 0.0 27.36 179.36 29.07 ;
   RECT 0.0 29.07 179.36 30.78 ;
   RECT 0.0 30.78 179.36 32.49 ;
   RECT 0.0 32.49 179.36 34.2 ;
   RECT 0.0 34.2 179.36 35.91 ;
   RECT 0.0 35.91 179.36 37.62 ;
   RECT 0.0 37.62 179.36 39.33 ;
   RECT 0.0 39.33 179.36 41.04 ;
   RECT 0.0 41.04 179.36 42.75 ;
   RECT 0.0 42.75 179.36 44.46 ;
   RECT 0.0 44.46 179.36 46.17 ;
   RECT 0.0 46.17 179.36 47.88 ;
   RECT 0.0 47.88 179.36 49.59 ;
   RECT 0.0 49.59 179.36 51.3 ;
   RECT 0.0 51.3 179.36 53.01 ;
   RECT 0.0 53.01 179.36 54.72 ;
   RECT 0.0 54.72 179.36 56.43 ;
   RECT 0.0 56.43 179.36 58.14 ;
   RECT 0.0 58.14 179.36 59.85 ;
   RECT 0.0 59.85 179.36 61.56 ;
   RECT 0.0 61.56 179.36 63.27 ;
   RECT 0.0 63.27 179.36 64.98 ;
   RECT 0.0 64.98 179.36 66.69 ;
   RECT 0.0 66.69 179.36 68.4 ;
   RECT 0.0 68.4 179.36 70.11 ;
   RECT 0.0 70.11 179.36 71.82 ;
   RECT 0.0 71.82 179.36 73.53 ;
   RECT 0.0 73.53 179.36 75.24 ;
   RECT 0.0 75.24 179.36 76.95 ;
   RECT 0.0 76.95 179.36 78.66 ;
   RECT 0.0 78.66 179.36 80.37 ;
   RECT 0.0 80.37 179.36 82.08 ;
   RECT 0.0 82.08 179.36 83.79 ;
   RECT 0.0 83.79 179.36 85.5 ;
   RECT 0.0 85.5 179.36 87.21 ;
   RECT 0.0 87.21 179.36 88.92 ;
   RECT 0.0 88.92 179.36 90.63 ;
   RECT 0.0 90.63 179.36 92.34 ;
   RECT 0.0 92.34 179.36 94.05 ;
   RECT 0.0 94.05 179.36 95.76 ;
   RECT 0.0 95.76 179.36 97.47 ;
   RECT 0.0 97.47 179.36 99.18 ;
   RECT 0.0 99.18 179.36 100.89 ;
   RECT 0.0 100.89 202.54 102.6 ;
   RECT 0.0 102.6 202.54 104.31 ;
   RECT 0.0 104.31 202.54 106.02 ;
   RECT 0.0 106.02 202.54 107.73 ;
   RECT 0.0 107.73 202.54 109.44 ;
   RECT 0.0 109.44 202.54 111.15 ;
   RECT 0.0 111.15 202.54 112.86 ;
   RECT 0.0 112.86 202.54 114.57 ;
   RECT 0.0 114.57 202.54 116.28 ;
   RECT 0.0 116.28 202.54 117.99 ;
   RECT 0.0 117.99 202.54 119.7 ;
   RECT 0.0 119.7 202.54 121.41 ;
   RECT 0.0 121.41 202.54 123.12 ;
   RECT 0.0 123.12 202.54 124.83 ;
   RECT 0.0 124.83 202.54 126.54 ;
   RECT 0.0 126.54 202.54 128.25 ;
   RECT 0.0 128.25 202.54 129.96 ;
   RECT 0.0 129.96 179.36 131.67 ;
   RECT 0.0 131.67 179.36 133.38 ;
   RECT 0.0 133.38 179.36 135.09 ;
   RECT 0.0 135.09 179.36 136.8 ;
   RECT 0.0 136.8 179.36 138.51 ;
   RECT 0.0 138.51 179.36 140.22 ;
   RECT 0.0 140.22 179.36 141.93 ;
   RECT 0.0 141.93 179.36 143.64 ;
   RECT 0.0 143.64 179.36 145.35 ;
   RECT 0.0 145.35 179.36 147.06 ;
   RECT 0.0 147.06 179.36 148.77 ;
   RECT 0.0 148.77 179.36 150.48 ;
   RECT 0.0 150.48 179.36 152.19 ;
   RECT 0.0 152.19 179.36 153.9 ;
   RECT 0.0 153.9 179.36 155.61 ;
   RECT 0.0 155.61 179.36 157.32 ;
   RECT 0.0 157.32 179.36 159.03 ;
   RECT 0.0 159.03 179.36 160.74 ;
   RECT 0.0 160.74 179.36 162.45 ;
   RECT 0.0 162.45 179.36 164.16 ;
   RECT 0.0 164.16 179.36 165.87 ;
   RECT 0.0 165.87 179.36 167.58 ;
   RECT 0.0 167.58 179.36 169.29 ;
   RECT 0.0 169.29 179.36 171.0 ;
   RECT 0.0 171.0 179.36 172.71 ;
   RECT 0.0 172.71 179.36 174.42 ;
   RECT 0.0 174.42 179.36 176.13 ;
   RECT 0.0 176.13 179.36 177.84 ;
   RECT 0.0 177.84 179.36 179.55 ;
   RECT 0.0 179.55 179.36 181.26 ;
   RECT 0.0 181.26 179.36 182.97 ;
   RECT 0.0 182.97 179.36 184.68 ;
   RECT 0.0 184.68 179.36 186.39 ;
   RECT 0.0 186.39 179.36 188.1 ;
   RECT 0.0 188.1 179.36 189.81 ;
   RECT 0.0 189.81 179.36 191.52 ;
   RECT 0.0 191.52 179.36 193.23 ;
   RECT 0.0 193.23 179.36 194.94 ;
   RECT 0.0 194.94 179.36 196.65 ;
   RECT 0.0 196.65 179.36 198.36 ;
   RECT 0.0 198.36 179.36 200.07 ;
   RECT 0.0 200.07 179.36 201.78 ;
   RECT 0.0 201.78 179.36 203.49 ;
   RECT 0.0 203.49 179.36 205.2 ;
   RECT 0.0 205.2 179.36 206.91 ;
   RECT 0.0 206.91 179.36 208.62 ;
   RECT 0.0 208.62 179.36 210.33 ;
   RECT 0.0 210.33 179.36 212.04 ;
   RECT 0.0 212.04 179.36 213.75 ;
  LAYER via1 ;
   RECT 0.0 0.0 179.36 1.71 ;
   RECT 0.0 1.71 179.36 3.42 ;
   RECT 0.0 3.42 179.36 5.13 ;
   RECT 0.0 5.13 179.36 6.84 ;
   RECT 0.0 6.84 179.36 8.55 ;
   RECT 0.0 8.55 179.36 10.26 ;
   RECT 0.0 10.26 179.36 11.97 ;
   RECT 0.0 11.97 179.36 13.68 ;
   RECT 0.0 13.68 179.36 15.39 ;
   RECT 0.0 15.39 179.36 17.1 ;
   RECT 0.0 17.1 179.36 18.81 ;
   RECT 0.0 18.81 179.36 20.52 ;
   RECT 0.0 20.52 179.36 22.23 ;
   RECT 0.0 22.23 179.36 23.94 ;
   RECT 0.0 23.94 179.36 25.65 ;
   RECT 0.0 25.65 179.36 27.36 ;
   RECT 0.0 27.36 179.36 29.07 ;
   RECT 0.0 29.07 179.36 30.78 ;
   RECT 0.0 30.78 179.36 32.49 ;
   RECT 0.0 32.49 179.36 34.2 ;
   RECT 0.0 34.2 179.36 35.91 ;
   RECT 0.0 35.91 179.36 37.62 ;
   RECT 0.0 37.62 179.36 39.33 ;
   RECT 0.0 39.33 179.36 41.04 ;
   RECT 0.0 41.04 179.36 42.75 ;
   RECT 0.0 42.75 179.36 44.46 ;
   RECT 0.0 44.46 179.36 46.17 ;
   RECT 0.0 46.17 179.36 47.88 ;
   RECT 0.0 47.88 179.36 49.59 ;
   RECT 0.0 49.59 179.36 51.3 ;
   RECT 0.0 51.3 179.36 53.01 ;
   RECT 0.0 53.01 179.36 54.72 ;
   RECT 0.0 54.72 179.36 56.43 ;
   RECT 0.0 56.43 179.36 58.14 ;
   RECT 0.0 58.14 179.36 59.85 ;
   RECT 0.0 59.85 179.36 61.56 ;
   RECT 0.0 61.56 179.36 63.27 ;
   RECT 0.0 63.27 179.36 64.98 ;
   RECT 0.0 64.98 179.36 66.69 ;
   RECT 0.0 66.69 179.36 68.4 ;
   RECT 0.0 68.4 179.36 70.11 ;
   RECT 0.0 70.11 179.36 71.82 ;
   RECT 0.0 71.82 179.36 73.53 ;
   RECT 0.0 73.53 179.36 75.24 ;
   RECT 0.0 75.24 179.36 76.95 ;
   RECT 0.0 76.95 179.36 78.66 ;
   RECT 0.0 78.66 179.36 80.37 ;
   RECT 0.0 80.37 179.36 82.08 ;
   RECT 0.0 82.08 179.36 83.79 ;
   RECT 0.0 83.79 179.36 85.5 ;
   RECT 0.0 85.5 179.36 87.21 ;
   RECT 0.0 87.21 179.36 88.92 ;
   RECT 0.0 88.92 179.36 90.63 ;
   RECT 0.0 90.63 179.36 92.34 ;
   RECT 0.0 92.34 179.36 94.05 ;
   RECT 0.0 94.05 179.36 95.76 ;
   RECT 0.0 95.76 179.36 97.47 ;
   RECT 0.0 97.47 179.36 99.18 ;
   RECT 0.0 99.18 179.36 100.89 ;
   RECT 0.0 100.89 202.54 102.6 ;
   RECT 0.0 102.6 202.54 104.31 ;
   RECT 0.0 104.31 202.54 106.02 ;
   RECT 0.0 106.02 202.54 107.73 ;
   RECT 0.0 107.73 202.54 109.44 ;
   RECT 0.0 109.44 202.54 111.15 ;
   RECT 0.0 111.15 202.54 112.86 ;
   RECT 0.0 112.86 202.54 114.57 ;
   RECT 0.0 114.57 202.54 116.28 ;
   RECT 0.0 116.28 202.54 117.99 ;
   RECT 0.0 117.99 202.54 119.7 ;
   RECT 0.0 119.7 202.54 121.41 ;
   RECT 0.0 121.41 202.54 123.12 ;
   RECT 0.0 123.12 202.54 124.83 ;
   RECT 0.0 124.83 202.54 126.54 ;
   RECT 0.0 126.54 202.54 128.25 ;
   RECT 0.0 128.25 202.54 129.96 ;
   RECT 0.0 129.96 179.36 131.67 ;
   RECT 0.0 131.67 179.36 133.38 ;
   RECT 0.0 133.38 179.36 135.09 ;
   RECT 0.0 135.09 179.36 136.8 ;
   RECT 0.0 136.8 179.36 138.51 ;
   RECT 0.0 138.51 179.36 140.22 ;
   RECT 0.0 140.22 179.36 141.93 ;
   RECT 0.0 141.93 179.36 143.64 ;
   RECT 0.0 143.64 179.36 145.35 ;
   RECT 0.0 145.35 179.36 147.06 ;
   RECT 0.0 147.06 179.36 148.77 ;
   RECT 0.0 148.77 179.36 150.48 ;
   RECT 0.0 150.48 179.36 152.19 ;
   RECT 0.0 152.19 179.36 153.9 ;
   RECT 0.0 153.9 179.36 155.61 ;
   RECT 0.0 155.61 179.36 157.32 ;
   RECT 0.0 157.32 179.36 159.03 ;
   RECT 0.0 159.03 179.36 160.74 ;
   RECT 0.0 160.74 179.36 162.45 ;
   RECT 0.0 162.45 179.36 164.16 ;
   RECT 0.0 164.16 179.36 165.87 ;
   RECT 0.0 165.87 179.36 167.58 ;
   RECT 0.0 167.58 179.36 169.29 ;
   RECT 0.0 169.29 179.36 171.0 ;
   RECT 0.0 171.0 179.36 172.71 ;
   RECT 0.0 172.71 179.36 174.42 ;
   RECT 0.0 174.42 179.36 176.13 ;
   RECT 0.0 176.13 179.36 177.84 ;
   RECT 0.0 177.84 179.36 179.55 ;
   RECT 0.0 179.55 179.36 181.26 ;
   RECT 0.0 181.26 179.36 182.97 ;
   RECT 0.0 182.97 179.36 184.68 ;
   RECT 0.0 184.68 179.36 186.39 ;
   RECT 0.0 186.39 179.36 188.1 ;
   RECT 0.0 188.1 179.36 189.81 ;
   RECT 0.0 189.81 179.36 191.52 ;
   RECT 0.0 191.52 179.36 193.23 ;
   RECT 0.0 193.23 179.36 194.94 ;
   RECT 0.0 194.94 179.36 196.65 ;
   RECT 0.0 196.65 179.36 198.36 ;
   RECT 0.0 198.36 179.36 200.07 ;
   RECT 0.0 200.07 179.36 201.78 ;
   RECT 0.0 201.78 179.36 203.49 ;
   RECT 0.0 203.49 179.36 205.2 ;
   RECT 0.0 205.2 179.36 206.91 ;
   RECT 0.0 206.91 179.36 208.62 ;
   RECT 0.0 208.62 179.36 210.33 ;
   RECT 0.0 210.33 179.36 212.04 ;
   RECT 0.0 212.04 179.36 213.75 ;
  LAYER metal2 ;
   RECT 0.0 0.0 179.36 1.71 ;
   RECT 0.0 1.71 179.36 3.42 ;
   RECT 0.0 3.42 179.36 5.13 ;
   RECT 0.0 5.13 179.36 6.84 ;
   RECT 0.0 6.84 179.36 8.55 ;
   RECT 0.0 8.55 179.36 10.26 ;
   RECT 0.0 10.26 179.36 11.97 ;
   RECT 0.0 11.97 179.36 13.68 ;
   RECT 0.0 13.68 179.36 15.39 ;
   RECT 0.0 15.39 179.36 17.1 ;
   RECT 0.0 17.1 179.36 18.81 ;
   RECT 0.0 18.81 179.36 20.52 ;
   RECT 0.0 20.52 179.36 22.23 ;
   RECT 0.0 22.23 179.36 23.94 ;
   RECT 0.0 23.94 179.36 25.65 ;
   RECT 0.0 25.65 179.36 27.36 ;
   RECT 0.0 27.36 179.36 29.07 ;
   RECT 0.0 29.07 179.36 30.78 ;
   RECT 0.0 30.78 179.36 32.49 ;
   RECT 0.0 32.49 179.36 34.2 ;
   RECT 0.0 34.2 179.36 35.91 ;
   RECT 0.0 35.91 179.36 37.62 ;
   RECT 0.0 37.62 179.36 39.33 ;
   RECT 0.0 39.33 179.36 41.04 ;
   RECT 0.0 41.04 179.36 42.75 ;
   RECT 0.0 42.75 179.36 44.46 ;
   RECT 0.0 44.46 179.36 46.17 ;
   RECT 0.0 46.17 179.36 47.88 ;
   RECT 0.0 47.88 179.36 49.59 ;
   RECT 0.0 49.59 179.36 51.3 ;
   RECT 0.0 51.3 179.36 53.01 ;
   RECT 0.0 53.01 179.36 54.72 ;
   RECT 0.0 54.72 179.36 56.43 ;
   RECT 0.0 56.43 179.36 58.14 ;
   RECT 0.0 58.14 179.36 59.85 ;
   RECT 0.0 59.85 179.36 61.56 ;
   RECT 0.0 61.56 179.36 63.27 ;
   RECT 0.0 63.27 179.36 64.98 ;
   RECT 0.0 64.98 179.36 66.69 ;
   RECT 0.0 66.69 179.36 68.4 ;
   RECT 0.0 68.4 179.36 70.11 ;
   RECT 0.0 70.11 179.36 71.82 ;
   RECT 0.0 71.82 179.36 73.53 ;
   RECT 0.0 73.53 179.36 75.24 ;
   RECT 0.0 75.24 179.36 76.95 ;
   RECT 0.0 76.95 179.36 78.66 ;
   RECT 0.0 78.66 179.36 80.37 ;
   RECT 0.0 80.37 179.36 82.08 ;
   RECT 0.0 82.08 179.36 83.79 ;
   RECT 0.0 83.79 179.36 85.5 ;
   RECT 0.0 85.5 179.36 87.21 ;
   RECT 0.0 87.21 179.36 88.92 ;
   RECT 0.0 88.92 179.36 90.63 ;
   RECT 0.0 90.63 179.36 92.34 ;
   RECT 0.0 92.34 179.36 94.05 ;
   RECT 0.0 94.05 179.36 95.76 ;
   RECT 0.0 95.76 179.36 97.47 ;
   RECT 0.0 97.47 179.36 99.18 ;
   RECT 0.0 99.18 179.36 100.89 ;
   RECT 0.0 100.89 202.54 102.6 ;
   RECT 0.0 102.6 202.54 104.31 ;
   RECT 0.0 104.31 202.54 106.02 ;
   RECT 0.0 106.02 202.54 107.73 ;
   RECT 0.0 107.73 202.54 109.44 ;
   RECT 0.0 109.44 202.54 111.15 ;
   RECT 0.0 111.15 202.54 112.86 ;
   RECT 0.0 112.86 202.54 114.57 ;
   RECT 0.0 114.57 202.54 116.28 ;
   RECT 0.0 116.28 202.54 117.99 ;
   RECT 0.0 117.99 202.54 119.7 ;
   RECT 0.0 119.7 202.54 121.41 ;
   RECT 0.0 121.41 202.54 123.12 ;
   RECT 0.0 123.12 202.54 124.83 ;
   RECT 0.0 124.83 202.54 126.54 ;
   RECT 0.0 126.54 202.54 128.25 ;
   RECT 0.0 128.25 202.54 129.96 ;
   RECT 0.0 129.96 179.36 131.67 ;
   RECT 0.0 131.67 179.36 133.38 ;
   RECT 0.0 133.38 179.36 135.09 ;
   RECT 0.0 135.09 179.36 136.8 ;
   RECT 0.0 136.8 179.36 138.51 ;
   RECT 0.0 138.51 179.36 140.22 ;
   RECT 0.0 140.22 179.36 141.93 ;
   RECT 0.0 141.93 179.36 143.64 ;
   RECT 0.0 143.64 179.36 145.35 ;
   RECT 0.0 145.35 179.36 147.06 ;
   RECT 0.0 147.06 179.36 148.77 ;
   RECT 0.0 148.77 179.36 150.48 ;
   RECT 0.0 150.48 179.36 152.19 ;
   RECT 0.0 152.19 179.36 153.9 ;
   RECT 0.0 153.9 179.36 155.61 ;
   RECT 0.0 155.61 179.36 157.32 ;
   RECT 0.0 157.32 179.36 159.03 ;
   RECT 0.0 159.03 179.36 160.74 ;
   RECT 0.0 160.74 179.36 162.45 ;
   RECT 0.0 162.45 179.36 164.16 ;
   RECT 0.0 164.16 179.36 165.87 ;
   RECT 0.0 165.87 179.36 167.58 ;
   RECT 0.0 167.58 179.36 169.29 ;
   RECT 0.0 169.29 179.36 171.0 ;
   RECT 0.0 171.0 179.36 172.71 ;
   RECT 0.0 172.71 179.36 174.42 ;
   RECT 0.0 174.42 179.36 176.13 ;
   RECT 0.0 176.13 179.36 177.84 ;
   RECT 0.0 177.84 179.36 179.55 ;
   RECT 0.0 179.55 179.36 181.26 ;
   RECT 0.0 181.26 179.36 182.97 ;
   RECT 0.0 182.97 179.36 184.68 ;
   RECT 0.0 184.68 179.36 186.39 ;
   RECT 0.0 186.39 179.36 188.1 ;
   RECT 0.0 188.1 179.36 189.81 ;
   RECT 0.0 189.81 179.36 191.52 ;
   RECT 0.0 191.52 179.36 193.23 ;
   RECT 0.0 193.23 179.36 194.94 ;
   RECT 0.0 194.94 179.36 196.65 ;
   RECT 0.0 196.65 179.36 198.36 ;
   RECT 0.0 198.36 179.36 200.07 ;
   RECT 0.0 200.07 179.36 201.78 ;
   RECT 0.0 201.78 179.36 203.49 ;
   RECT 0.0 203.49 179.36 205.2 ;
   RECT 0.0 205.2 179.36 206.91 ;
   RECT 0.0 206.91 179.36 208.62 ;
   RECT 0.0 208.62 179.36 210.33 ;
   RECT 0.0 210.33 179.36 212.04 ;
   RECT 0.0 212.04 179.36 213.75 ;
  LAYER via2 ;
   RECT 0.0 0.0 179.36 1.71 ;
   RECT 0.0 1.71 179.36 3.42 ;
   RECT 0.0 3.42 179.36 5.13 ;
   RECT 0.0 5.13 179.36 6.84 ;
   RECT 0.0 6.84 179.36 8.55 ;
   RECT 0.0 8.55 179.36 10.26 ;
   RECT 0.0 10.26 179.36 11.97 ;
   RECT 0.0 11.97 179.36 13.68 ;
   RECT 0.0 13.68 179.36 15.39 ;
   RECT 0.0 15.39 179.36 17.1 ;
   RECT 0.0 17.1 179.36 18.81 ;
   RECT 0.0 18.81 179.36 20.52 ;
   RECT 0.0 20.52 179.36 22.23 ;
   RECT 0.0 22.23 179.36 23.94 ;
   RECT 0.0 23.94 179.36 25.65 ;
   RECT 0.0 25.65 179.36 27.36 ;
   RECT 0.0 27.36 179.36 29.07 ;
   RECT 0.0 29.07 179.36 30.78 ;
   RECT 0.0 30.78 179.36 32.49 ;
   RECT 0.0 32.49 179.36 34.2 ;
   RECT 0.0 34.2 179.36 35.91 ;
   RECT 0.0 35.91 179.36 37.62 ;
   RECT 0.0 37.62 179.36 39.33 ;
   RECT 0.0 39.33 179.36 41.04 ;
   RECT 0.0 41.04 179.36 42.75 ;
   RECT 0.0 42.75 179.36 44.46 ;
   RECT 0.0 44.46 179.36 46.17 ;
   RECT 0.0 46.17 179.36 47.88 ;
   RECT 0.0 47.88 179.36 49.59 ;
   RECT 0.0 49.59 179.36 51.3 ;
   RECT 0.0 51.3 179.36 53.01 ;
   RECT 0.0 53.01 179.36 54.72 ;
   RECT 0.0 54.72 179.36 56.43 ;
   RECT 0.0 56.43 179.36 58.14 ;
   RECT 0.0 58.14 179.36 59.85 ;
   RECT 0.0 59.85 179.36 61.56 ;
   RECT 0.0 61.56 179.36 63.27 ;
   RECT 0.0 63.27 179.36 64.98 ;
   RECT 0.0 64.98 179.36 66.69 ;
   RECT 0.0 66.69 179.36 68.4 ;
   RECT 0.0 68.4 179.36 70.11 ;
   RECT 0.0 70.11 179.36 71.82 ;
   RECT 0.0 71.82 179.36 73.53 ;
   RECT 0.0 73.53 179.36 75.24 ;
   RECT 0.0 75.24 179.36 76.95 ;
   RECT 0.0 76.95 179.36 78.66 ;
   RECT 0.0 78.66 179.36 80.37 ;
   RECT 0.0 80.37 179.36 82.08 ;
   RECT 0.0 82.08 179.36 83.79 ;
   RECT 0.0 83.79 179.36 85.5 ;
   RECT 0.0 85.5 179.36 87.21 ;
   RECT 0.0 87.21 179.36 88.92 ;
   RECT 0.0 88.92 179.36 90.63 ;
   RECT 0.0 90.63 179.36 92.34 ;
   RECT 0.0 92.34 179.36 94.05 ;
   RECT 0.0 94.05 179.36 95.76 ;
   RECT 0.0 95.76 179.36 97.47 ;
   RECT 0.0 97.47 179.36 99.18 ;
   RECT 0.0 99.18 179.36 100.89 ;
   RECT 0.0 100.89 202.54 102.6 ;
   RECT 0.0 102.6 202.54 104.31 ;
   RECT 0.0 104.31 202.54 106.02 ;
   RECT 0.0 106.02 202.54 107.73 ;
   RECT 0.0 107.73 202.54 109.44 ;
   RECT 0.0 109.44 202.54 111.15 ;
   RECT 0.0 111.15 202.54 112.86 ;
   RECT 0.0 112.86 202.54 114.57 ;
   RECT 0.0 114.57 202.54 116.28 ;
   RECT 0.0 116.28 202.54 117.99 ;
   RECT 0.0 117.99 202.54 119.7 ;
   RECT 0.0 119.7 202.54 121.41 ;
   RECT 0.0 121.41 202.54 123.12 ;
   RECT 0.0 123.12 202.54 124.83 ;
   RECT 0.0 124.83 202.54 126.54 ;
   RECT 0.0 126.54 202.54 128.25 ;
   RECT 0.0 128.25 202.54 129.96 ;
   RECT 0.0 129.96 179.36 131.67 ;
   RECT 0.0 131.67 179.36 133.38 ;
   RECT 0.0 133.38 179.36 135.09 ;
   RECT 0.0 135.09 179.36 136.8 ;
   RECT 0.0 136.8 179.36 138.51 ;
   RECT 0.0 138.51 179.36 140.22 ;
   RECT 0.0 140.22 179.36 141.93 ;
   RECT 0.0 141.93 179.36 143.64 ;
   RECT 0.0 143.64 179.36 145.35 ;
   RECT 0.0 145.35 179.36 147.06 ;
   RECT 0.0 147.06 179.36 148.77 ;
   RECT 0.0 148.77 179.36 150.48 ;
   RECT 0.0 150.48 179.36 152.19 ;
   RECT 0.0 152.19 179.36 153.9 ;
   RECT 0.0 153.9 179.36 155.61 ;
   RECT 0.0 155.61 179.36 157.32 ;
   RECT 0.0 157.32 179.36 159.03 ;
   RECT 0.0 159.03 179.36 160.74 ;
   RECT 0.0 160.74 179.36 162.45 ;
   RECT 0.0 162.45 179.36 164.16 ;
   RECT 0.0 164.16 179.36 165.87 ;
   RECT 0.0 165.87 179.36 167.58 ;
   RECT 0.0 167.58 179.36 169.29 ;
   RECT 0.0 169.29 179.36 171.0 ;
   RECT 0.0 171.0 179.36 172.71 ;
   RECT 0.0 172.71 179.36 174.42 ;
   RECT 0.0 174.42 179.36 176.13 ;
   RECT 0.0 176.13 179.36 177.84 ;
   RECT 0.0 177.84 179.36 179.55 ;
   RECT 0.0 179.55 179.36 181.26 ;
   RECT 0.0 181.26 179.36 182.97 ;
   RECT 0.0 182.97 179.36 184.68 ;
   RECT 0.0 184.68 179.36 186.39 ;
   RECT 0.0 186.39 179.36 188.1 ;
   RECT 0.0 188.1 179.36 189.81 ;
   RECT 0.0 189.81 179.36 191.52 ;
   RECT 0.0 191.52 179.36 193.23 ;
   RECT 0.0 193.23 179.36 194.94 ;
   RECT 0.0 194.94 179.36 196.65 ;
   RECT 0.0 196.65 179.36 198.36 ;
   RECT 0.0 198.36 179.36 200.07 ;
   RECT 0.0 200.07 179.36 201.78 ;
   RECT 0.0 201.78 179.36 203.49 ;
   RECT 0.0 203.49 179.36 205.2 ;
   RECT 0.0 205.2 179.36 206.91 ;
   RECT 0.0 206.91 179.36 208.62 ;
   RECT 0.0 208.62 179.36 210.33 ;
   RECT 0.0 210.33 179.36 212.04 ;
   RECT 0.0 212.04 179.36 213.75 ;
  LAYER metal3 ;
   RECT 0.0 0.0 179.36 1.71 ;
   RECT 0.0 1.71 179.36 3.42 ;
   RECT 0.0 3.42 179.36 5.13 ;
   RECT 0.0 5.13 179.36 6.84 ;
   RECT 0.0 6.84 179.36 8.55 ;
   RECT 0.0 8.55 179.36 10.26 ;
   RECT 0.0 10.26 179.36 11.97 ;
   RECT 0.0 11.97 179.36 13.68 ;
   RECT 0.0 13.68 179.36 15.39 ;
   RECT 0.0 15.39 179.36 17.1 ;
   RECT 0.0 17.1 179.36 18.81 ;
   RECT 0.0 18.81 179.36 20.52 ;
   RECT 0.0 20.52 179.36 22.23 ;
   RECT 0.0 22.23 179.36 23.94 ;
   RECT 0.0 23.94 179.36 25.65 ;
   RECT 0.0 25.65 179.36 27.36 ;
   RECT 0.0 27.36 179.36 29.07 ;
   RECT 0.0 29.07 179.36 30.78 ;
   RECT 0.0 30.78 179.36 32.49 ;
   RECT 0.0 32.49 179.36 34.2 ;
   RECT 0.0 34.2 179.36 35.91 ;
   RECT 0.0 35.91 179.36 37.62 ;
   RECT 0.0 37.62 179.36 39.33 ;
   RECT 0.0 39.33 179.36 41.04 ;
   RECT 0.0 41.04 179.36 42.75 ;
   RECT 0.0 42.75 179.36 44.46 ;
   RECT 0.0 44.46 179.36 46.17 ;
   RECT 0.0 46.17 179.36 47.88 ;
   RECT 0.0 47.88 179.36 49.59 ;
   RECT 0.0 49.59 179.36 51.3 ;
   RECT 0.0 51.3 179.36 53.01 ;
   RECT 0.0 53.01 179.36 54.72 ;
   RECT 0.0 54.72 179.36 56.43 ;
   RECT 0.0 56.43 179.36 58.14 ;
   RECT 0.0 58.14 179.36 59.85 ;
   RECT 0.0 59.85 179.36 61.56 ;
   RECT 0.0 61.56 179.36 63.27 ;
   RECT 0.0 63.27 179.36 64.98 ;
   RECT 0.0 64.98 179.36 66.69 ;
   RECT 0.0 66.69 179.36 68.4 ;
   RECT 0.0 68.4 179.36 70.11 ;
   RECT 0.0 70.11 179.36 71.82 ;
   RECT 0.0 71.82 179.36 73.53 ;
   RECT 0.0 73.53 179.36 75.24 ;
   RECT 0.0 75.24 179.36 76.95 ;
   RECT 0.0 76.95 179.36 78.66 ;
   RECT 0.0 78.66 179.36 80.37 ;
   RECT 0.0 80.37 179.36 82.08 ;
   RECT 0.0 82.08 179.36 83.79 ;
   RECT 0.0 83.79 179.36 85.5 ;
   RECT 0.0 85.5 179.36 87.21 ;
   RECT 0.0 87.21 179.36 88.92 ;
   RECT 0.0 88.92 179.36 90.63 ;
   RECT 0.0 90.63 179.36 92.34 ;
   RECT 0.0 92.34 179.36 94.05 ;
   RECT 0.0 94.05 179.36 95.76 ;
   RECT 0.0 95.76 179.36 97.47 ;
   RECT 0.0 97.47 179.36 99.18 ;
   RECT 0.0 99.18 179.36 100.89 ;
   RECT 0.0 100.89 202.54 102.6 ;
   RECT 0.0 102.6 202.54 104.31 ;
   RECT 0.0 104.31 202.54 106.02 ;
   RECT 0.0 106.02 202.54 107.73 ;
   RECT 0.0 107.73 202.54 109.44 ;
   RECT 0.0 109.44 202.54 111.15 ;
   RECT 0.0 111.15 202.54 112.86 ;
   RECT 0.0 112.86 202.54 114.57 ;
   RECT 0.0 114.57 202.54 116.28 ;
   RECT 0.0 116.28 202.54 117.99 ;
   RECT 0.0 117.99 202.54 119.7 ;
   RECT 0.0 119.7 202.54 121.41 ;
   RECT 0.0 121.41 202.54 123.12 ;
   RECT 0.0 123.12 202.54 124.83 ;
   RECT 0.0 124.83 202.54 126.54 ;
   RECT 0.0 126.54 202.54 128.25 ;
   RECT 0.0 128.25 202.54 129.96 ;
   RECT 0.0 129.96 179.36 131.67 ;
   RECT 0.0 131.67 179.36 133.38 ;
   RECT 0.0 133.38 179.36 135.09 ;
   RECT 0.0 135.09 179.36 136.8 ;
   RECT 0.0 136.8 179.36 138.51 ;
   RECT 0.0 138.51 179.36 140.22 ;
   RECT 0.0 140.22 179.36 141.93 ;
   RECT 0.0 141.93 179.36 143.64 ;
   RECT 0.0 143.64 179.36 145.35 ;
   RECT 0.0 145.35 179.36 147.06 ;
   RECT 0.0 147.06 179.36 148.77 ;
   RECT 0.0 148.77 179.36 150.48 ;
   RECT 0.0 150.48 179.36 152.19 ;
   RECT 0.0 152.19 179.36 153.9 ;
   RECT 0.0 153.9 179.36 155.61 ;
   RECT 0.0 155.61 179.36 157.32 ;
   RECT 0.0 157.32 179.36 159.03 ;
   RECT 0.0 159.03 179.36 160.74 ;
   RECT 0.0 160.74 179.36 162.45 ;
   RECT 0.0 162.45 179.36 164.16 ;
   RECT 0.0 164.16 179.36 165.87 ;
   RECT 0.0 165.87 179.36 167.58 ;
   RECT 0.0 167.58 179.36 169.29 ;
   RECT 0.0 169.29 179.36 171.0 ;
   RECT 0.0 171.0 179.36 172.71 ;
   RECT 0.0 172.71 179.36 174.42 ;
   RECT 0.0 174.42 179.36 176.13 ;
   RECT 0.0 176.13 179.36 177.84 ;
   RECT 0.0 177.84 179.36 179.55 ;
   RECT 0.0 179.55 179.36 181.26 ;
   RECT 0.0 181.26 179.36 182.97 ;
   RECT 0.0 182.97 179.36 184.68 ;
   RECT 0.0 184.68 179.36 186.39 ;
   RECT 0.0 186.39 179.36 188.1 ;
   RECT 0.0 188.1 179.36 189.81 ;
   RECT 0.0 189.81 179.36 191.52 ;
   RECT 0.0 191.52 179.36 193.23 ;
   RECT 0.0 193.23 179.36 194.94 ;
   RECT 0.0 194.94 179.36 196.65 ;
   RECT 0.0 196.65 179.36 198.36 ;
   RECT 0.0 198.36 179.36 200.07 ;
   RECT 0.0 200.07 179.36 201.78 ;
   RECT 0.0 201.78 179.36 203.49 ;
   RECT 0.0 203.49 179.36 205.2 ;
   RECT 0.0 205.2 179.36 206.91 ;
   RECT 0.0 206.91 179.36 208.62 ;
   RECT 0.0 208.62 179.36 210.33 ;
   RECT 0.0 210.33 179.36 212.04 ;
   RECT 0.0 212.04 179.36 213.75 ;
  LAYER via3 ;
   RECT 0.0 0.0 179.36 1.71 ;
   RECT 0.0 1.71 179.36 3.42 ;
   RECT 0.0 3.42 179.36 5.13 ;
   RECT 0.0 5.13 179.36 6.84 ;
   RECT 0.0 6.84 179.36 8.55 ;
   RECT 0.0 8.55 179.36 10.26 ;
   RECT 0.0 10.26 179.36 11.97 ;
   RECT 0.0 11.97 179.36 13.68 ;
   RECT 0.0 13.68 179.36 15.39 ;
   RECT 0.0 15.39 179.36 17.1 ;
   RECT 0.0 17.1 179.36 18.81 ;
   RECT 0.0 18.81 179.36 20.52 ;
   RECT 0.0 20.52 179.36 22.23 ;
   RECT 0.0 22.23 179.36 23.94 ;
   RECT 0.0 23.94 179.36 25.65 ;
   RECT 0.0 25.65 179.36 27.36 ;
   RECT 0.0 27.36 179.36 29.07 ;
   RECT 0.0 29.07 179.36 30.78 ;
   RECT 0.0 30.78 179.36 32.49 ;
   RECT 0.0 32.49 179.36 34.2 ;
   RECT 0.0 34.2 179.36 35.91 ;
   RECT 0.0 35.91 179.36 37.62 ;
   RECT 0.0 37.62 179.36 39.33 ;
   RECT 0.0 39.33 179.36 41.04 ;
   RECT 0.0 41.04 179.36 42.75 ;
   RECT 0.0 42.75 179.36 44.46 ;
   RECT 0.0 44.46 179.36 46.17 ;
   RECT 0.0 46.17 179.36 47.88 ;
   RECT 0.0 47.88 179.36 49.59 ;
   RECT 0.0 49.59 179.36 51.3 ;
   RECT 0.0 51.3 179.36 53.01 ;
   RECT 0.0 53.01 179.36 54.72 ;
   RECT 0.0 54.72 179.36 56.43 ;
   RECT 0.0 56.43 179.36 58.14 ;
   RECT 0.0 58.14 179.36 59.85 ;
   RECT 0.0 59.85 179.36 61.56 ;
   RECT 0.0 61.56 179.36 63.27 ;
   RECT 0.0 63.27 179.36 64.98 ;
   RECT 0.0 64.98 179.36 66.69 ;
   RECT 0.0 66.69 179.36 68.4 ;
   RECT 0.0 68.4 179.36 70.11 ;
   RECT 0.0 70.11 179.36 71.82 ;
   RECT 0.0 71.82 179.36 73.53 ;
   RECT 0.0 73.53 179.36 75.24 ;
   RECT 0.0 75.24 179.36 76.95 ;
   RECT 0.0 76.95 179.36 78.66 ;
   RECT 0.0 78.66 179.36 80.37 ;
   RECT 0.0 80.37 179.36 82.08 ;
   RECT 0.0 82.08 179.36 83.79 ;
   RECT 0.0 83.79 179.36 85.5 ;
   RECT 0.0 85.5 179.36 87.21 ;
   RECT 0.0 87.21 179.36 88.92 ;
   RECT 0.0 88.92 179.36 90.63 ;
   RECT 0.0 90.63 179.36 92.34 ;
   RECT 0.0 92.34 179.36 94.05 ;
   RECT 0.0 94.05 179.36 95.76 ;
   RECT 0.0 95.76 179.36 97.47 ;
   RECT 0.0 97.47 179.36 99.18 ;
   RECT 0.0 99.18 179.36 100.89 ;
   RECT 0.0 100.89 202.54 102.6 ;
   RECT 0.0 102.6 202.54 104.31 ;
   RECT 0.0 104.31 202.54 106.02 ;
   RECT 0.0 106.02 202.54 107.73 ;
   RECT 0.0 107.73 202.54 109.44 ;
   RECT 0.0 109.44 202.54 111.15 ;
   RECT 0.0 111.15 202.54 112.86 ;
   RECT 0.0 112.86 202.54 114.57 ;
   RECT 0.0 114.57 202.54 116.28 ;
   RECT 0.0 116.28 202.54 117.99 ;
   RECT 0.0 117.99 202.54 119.7 ;
   RECT 0.0 119.7 202.54 121.41 ;
   RECT 0.0 121.41 202.54 123.12 ;
   RECT 0.0 123.12 202.54 124.83 ;
   RECT 0.0 124.83 202.54 126.54 ;
   RECT 0.0 126.54 202.54 128.25 ;
   RECT 0.0 128.25 202.54 129.96 ;
   RECT 0.0 129.96 179.36 131.67 ;
   RECT 0.0 131.67 179.36 133.38 ;
   RECT 0.0 133.38 179.36 135.09 ;
   RECT 0.0 135.09 179.36 136.8 ;
   RECT 0.0 136.8 179.36 138.51 ;
   RECT 0.0 138.51 179.36 140.22 ;
   RECT 0.0 140.22 179.36 141.93 ;
   RECT 0.0 141.93 179.36 143.64 ;
   RECT 0.0 143.64 179.36 145.35 ;
   RECT 0.0 145.35 179.36 147.06 ;
   RECT 0.0 147.06 179.36 148.77 ;
   RECT 0.0 148.77 179.36 150.48 ;
   RECT 0.0 150.48 179.36 152.19 ;
   RECT 0.0 152.19 179.36 153.9 ;
   RECT 0.0 153.9 179.36 155.61 ;
   RECT 0.0 155.61 179.36 157.32 ;
   RECT 0.0 157.32 179.36 159.03 ;
   RECT 0.0 159.03 179.36 160.74 ;
   RECT 0.0 160.74 179.36 162.45 ;
   RECT 0.0 162.45 179.36 164.16 ;
   RECT 0.0 164.16 179.36 165.87 ;
   RECT 0.0 165.87 179.36 167.58 ;
   RECT 0.0 167.58 179.36 169.29 ;
   RECT 0.0 169.29 179.36 171.0 ;
   RECT 0.0 171.0 179.36 172.71 ;
   RECT 0.0 172.71 179.36 174.42 ;
   RECT 0.0 174.42 179.36 176.13 ;
   RECT 0.0 176.13 179.36 177.84 ;
   RECT 0.0 177.84 179.36 179.55 ;
   RECT 0.0 179.55 179.36 181.26 ;
   RECT 0.0 181.26 179.36 182.97 ;
   RECT 0.0 182.97 179.36 184.68 ;
   RECT 0.0 184.68 179.36 186.39 ;
   RECT 0.0 186.39 179.36 188.1 ;
   RECT 0.0 188.1 179.36 189.81 ;
   RECT 0.0 189.81 179.36 191.52 ;
   RECT 0.0 191.52 179.36 193.23 ;
   RECT 0.0 193.23 179.36 194.94 ;
   RECT 0.0 194.94 179.36 196.65 ;
   RECT 0.0 196.65 179.36 198.36 ;
   RECT 0.0 198.36 179.36 200.07 ;
   RECT 0.0 200.07 179.36 201.78 ;
   RECT 0.0 201.78 179.36 203.49 ;
   RECT 0.0 203.49 179.36 205.2 ;
   RECT 0.0 205.2 179.36 206.91 ;
   RECT 0.0 206.91 179.36 208.62 ;
   RECT 0.0 208.62 179.36 210.33 ;
   RECT 0.0 210.33 179.36 212.04 ;
   RECT 0.0 212.04 179.36 213.75 ;
  LAYER metal4 ;
   RECT 0.0 0.0 179.36 1.71 ;
   RECT 0.0 1.71 179.36 3.42 ;
   RECT 0.0 3.42 179.36 5.13 ;
   RECT 0.0 5.13 179.36 6.84 ;
   RECT 0.0 6.84 179.36 8.55 ;
   RECT 0.0 8.55 179.36 10.26 ;
   RECT 0.0 10.26 179.36 11.97 ;
   RECT 0.0 11.97 179.36 13.68 ;
   RECT 0.0 13.68 179.36 15.39 ;
   RECT 0.0 15.39 179.36 17.1 ;
   RECT 0.0 17.1 179.36 18.81 ;
   RECT 0.0 18.81 179.36 20.52 ;
   RECT 0.0 20.52 179.36 22.23 ;
   RECT 0.0 22.23 179.36 23.94 ;
   RECT 0.0 23.94 179.36 25.65 ;
   RECT 0.0 25.65 179.36 27.36 ;
   RECT 0.0 27.36 179.36 29.07 ;
   RECT 0.0 29.07 179.36 30.78 ;
   RECT 0.0 30.78 179.36 32.49 ;
   RECT 0.0 32.49 179.36 34.2 ;
   RECT 0.0 34.2 179.36 35.91 ;
   RECT 0.0 35.91 179.36 37.62 ;
   RECT 0.0 37.62 179.36 39.33 ;
   RECT 0.0 39.33 179.36 41.04 ;
   RECT 0.0 41.04 179.36 42.75 ;
   RECT 0.0 42.75 179.36 44.46 ;
   RECT 0.0 44.46 179.36 46.17 ;
   RECT 0.0 46.17 179.36 47.88 ;
   RECT 0.0 47.88 179.36 49.59 ;
   RECT 0.0 49.59 179.36 51.3 ;
   RECT 0.0 51.3 179.36 53.01 ;
   RECT 0.0 53.01 179.36 54.72 ;
   RECT 0.0 54.72 179.36 56.43 ;
   RECT 0.0 56.43 179.36 58.14 ;
   RECT 0.0 58.14 179.36 59.85 ;
   RECT 0.0 59.85 179.36 61.56 ;
   RECT 0.0 61.56 179.36 63.27 ;
   RECT 0.0 63.27 179.36 64.98 ;
   RECT 0.0 64.98 179.36 66.69 ;
   RECT 0.0 66.69 179.36 68.4 ;
   RECT 0.0 68.4 179.36 70.11 ;
   RECT 0.0 70.11 179.36 71.82 ;
   RECT 0.0 71.82 179.36 73.53 ;
   RECT 0.0 73.53 179.36 75.24 ;
   RECT 0.0 75.24 179.36 76.95 ;
   RECT 0.0 76.95 179.36 78.66 ;
   RECT 0.0 78.66 179.36 80.37 ;
   RECT 0.0 80.37 179.36 82.08 ;
   RECT 0.0 82.08 179.36 83.79 ;
   RECT 0.0 83.79 179.36 85.5 ;
   RECT 0.0 85.5 179.36 87.21 ;
   RECT 0.0 87.21 179.36 88.92 ;
   RECT 0.0 88.92 179.36 90.63 ;
   RECT 0.0 90.63 179.36 92.34 ;
   RECT 0.0 92.34 179.36 94.05 ;
   RECT 0.0 94.05 179.36 95.76 ;
   RECT 0.0 95.76 179.36 97.47 ;
   RECT 0.0 97.47 179.36 99.18 ;
   RECT 0.0 99.18 179.36 100.89 ;
   RECT 0.0 100.89 202.54 102.6 ;
   RECT 0.0 102.6 202.54 104.31 ;
   RECT 0.0 104.31 202.54 106.02 ;
   RECT 0.0 106.02 202.54 107.73 ;
   RECT 0.0 107.73 202.54 109.44 ;
   RECT 0.0 109.44 202.54 111.15 ;
   RECT 0.0 111.15 202.54 112.86 ;
   RECT 0.0 112.86 202.54 114.57 ;
   RECT 0.0 114.57 202.54 116.28 ;
   RECT 0.0 116.28 202.54 117.99 ;
   RECT 0.0 117.99 202.54 119.7 ;
   RECT 0.0 119.7 202.54 121.41 ;
   RECT 0.0 121.41 202.54 123.12 ;
   RECT 0.0 123.12 202.54 124.83 ;
   RECT 0.0 124.83 202.54 126.54 ;
   RECT 0.0 126.54 202.54 128.25 ;
   RECT 0.0 128.25 202.54 129.96 ;
   RECT 0.0 129.96 179.36 131.67 ;
   RECT 0.0 131.67 179.36 133.38 ;
   RECT 0.0 133.38 179.36 135.09 ;
   RECT 0.0 135.09 179.36 136.8 ;
   RECT 0.0 136.8 179.36 138.51 ;
   RECT 0.0 138.51 179.36 140.22 ;
   RECT 0.0 140.22 179.36 141.93 ;
   RECT 0.0 141.93 179.36 143.64 ;
   RECT 0.0 143.64 179.36 145.35 ;
   RECT 0.0 145.35 179.36 147.06 ;
   RECT 0.0 147.06 179.36 148.77 ;
   RECT 0.0 148.77 179.36 150.48 ;
   RECT 0.0 150.48 179.36 152.19 ;
   RECT 0.0 152.19 179.36 153.9 ;
   RECT 0.0 153.9 179.36 155.61 ;
   RECT 0.0 155.61 179.36 157.32 ;
   RECT 0.0 157.32 179.36 159.03 ;
   RECT 0.0 159.03 179.36 160.74 ;
   RECT 0.0 160.74 179.36 162.45 ;
   RECT 0.0 162.45 179.36 164.16 ;
   RECT 0.0 164.16 179.36 165.87 ;
   RECT 0.0 165.87 179.36 167.58 ;
   RECT 0.0 167.58 179.36 169.29 ;
   RECT 0.0 169.29 179.36 171.0 ;
   RECT 0.0 171.0 179.36 172.71 ;
   RECT 0.0 172.71 179.36 174.42 ;
   RECT 0.0 174.42 179.36 176.13 ;
   RECT 0.0 176.13 179.36 177.84 ;
   RECT 0.0 177.84 179.36 179.55 ;
   RECT 0.0 179.55 179.36 181.26 ;
   RECT 0.0 181.26 179.36 182.97 ;
   RECT 0.0 182.97 179.36 184.68 ;
   RECT 0.0 184.68 179.36 186.39 ;
   RECT 0.0 186.39 179.36 188.1 ;
   RECT 0.0 188.1 179.36 189.81 ;
   RECT 0.0 189.81 179.36 191.52 ;
   RECT 0.0 191.52 179.36 193.23 ;
   RECT 0.0 193.23 179.36 194.94 ;
   RECT 0.0 194.94 179.36 196.65 ;
   RECT 0.0 196.65 179.36 198.36 ;
   RECT 0.0 198.36 179.36 200.07 ;
   RECT 0.0 200.07 179.36 201.78 ;
   RECT 0.0 201.78 179.36 203.49 ;
   RECT 0.0 203.49 179.36 205.2 ;
   RECT 0.0 205.2 179.36 206.91 ;
   RECT 0.0 206.91 179.36 208.62 ;
   RECT 0.0 208.62 179.36 210.33 ;
   RECT 0.0 210.33 179.36 212.04 ;
   RECT 0.0 212.04 179.36 213.75 ;
 END
END block_533x1125_87

MACRO block_341x369_74
 CLASS BLOCK ;
 FOREIGN block_341x369_74 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 129.58 BY 70.11 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 20.235 126.445 20.805 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 26.695 126.445 27.265 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 6.935 3.325 7.505 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 9.215 3.325 9.785 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 10.735 3.325 11.305 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 13.015 3.325 13.585 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 13.395 4.085 13.965 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 13.775 3.325 14.345 ;
  END
 END o7
 PIN o8
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 15.295 3.325 15.865 ;
  END
 END o8
 PIN o9
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 16.055 3.325 16.625 ;
  END
 END o9
 PIN o10
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 12.635 4.085 13.205 ;
  END
 END o10
 PIN o11
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 19.855 3.325 20.425 ;
  END
 END o11
 PIN o12
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 20.615 3.325 21.185 ;
  END
 END o12
 PIN o13
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 21.375 3.325 21.945 ;
  END
 END o13
 PIN o14
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 22.135 3.325 22.705 ;
  END
 END o14
 PIN o15
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 18.335 3.325 18.905 ;
  END
 END o15
 PIN o16
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 25.935 3.325 26.505 ;
  END
 END o16
 PIN o17
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 26.695 3.325 27.265 ;
  END
 END o17
 PIN o18
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 27.455 3.325 28.025 ;
  END
 END o18
 PIN o19
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 28.975 3.325 29.545 ;
  END
 END o19
 PIN o20
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 25.175 3.325 25.745 ;
  END
 END o20
 PIN o21
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 32.015 3.325 32.585 ;
  END
 END o21
 PIN o22
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 33.535 3.325 34.105 ;
  END
 END o22
 PIN o23
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 34.295 3.325 34.865 ;
  END
 END o23
 PIN o24
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 35.055 3.325 35.625 ;
  END
 END o24
 PIN o25
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 31.255 3.325 31.825 ;
  END
 END o25
 PIN o26
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 38.095 126.445 38.665 ;
  END
 END o26
 PIN o27
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 38.855 126.445 39.425 ;
  END
 END o27
 PIN o28
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 39.615 126.445 40.185 ;
  END
 END o28
 PIN o29
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 42.655 126.445 43.225 ;
  END
 END o29
 PIN o30
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 21.755 126.445 22.325 ;
  END
 END o30
 PIN o31
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 31.255 126.445 31.825 ;
  END
 END o31
 PIN o32
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 32.015 126.445 32.585 ;
  END
 END o32
 PIN o33
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 33.535 126.445 34.105 ;
  END
 END o33
 PIN o34
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 34.295 126.445 34.865 ;
  END
 END o34
 PIN o35
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 30.495 126.445 31.065 ;
  END
 END o35
 PIN o36
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 28.975 126.445 29.545 ;
  END
 END o36
 PIN o37
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 41.135 3.325 41.705 ;
  END
 END o37
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 35.815 126.445 36.385 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 43.035 125.685 43.605 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 32.395 125.685 32.965 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 35.435 125.685 36.005 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 36.955 126.445 37.525 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 36.575 125.685 37.145 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 33.915 125.685 34.485 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 30.115 125.685 30.685 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 40.375 3.325 40.945 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 8.455 3.325 9.025 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 25.935 126.445 26.505 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 25.175 126.445 25.745 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 24.415 126.445 24.985 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 34.675 125.685 35.245 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 30.875 125.685 31.445 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 40.755 126.445 41.325 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 27.455 126.445 28.025 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 38.475 125.685 39.045 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 39.995 125.685 40.565 ;
  END
 END i18
 PIN i19
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 39.235 125.685 39.805 ;
  END
 END i19
 PIN i20
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 124.355 40.375 124.925 40.945 ;
  END
 END i20
 PIN i21
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 8.455 126.445 9.025 ;
  END
 END i21
 PIN i22
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 9.215 126.445 9.785 ;
  END
 END i22
 PIN i23
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 10.735 126.445 11.305 ;
  END
 END i23
 PIN i24
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 11.495 126.445 12.065 ;
  END
 END i24
 PIN i25
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 12.255 126.445 12.825 ;
  END
 END i25
 PIN i26
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 13.015 126.445 13.585 ;
  END
 END i26
 PIN i27
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 8.075 125.685 8.645 ;
  END
 END i27
 PIN i28
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 7.695 126.445 8.265 ;
  END
 END i28
 PIN i29
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 7.315 125.685 7.885 ;
  END
 END i29
 PIN i30
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 6.935 126.445 7.505 ;
  END
 END i30
 PIN i31
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 6.555 125.685 7.125 ;
  END
 END i31
 PIN i32
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 13.775 126.445 14.345 ;
  END
 END i32
 PIN i33
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 15.295 126.445 15.865 ;
  END
 END i33
 PIN i34
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 16.055 126.445 16.625 ;
  END
 END i34
 PIN i35
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 16.815 126.445 17.385 ;
  END
 END i35
 OBS
  LAYER metal1 ;
   RECT 0 0 129.58 70.11 ;
  LAYER via1 ;
   RECT 0 0 129.58 70.11 ;
  LAYER metal2 ;
   RECT 0 0 129.58 70.11 ;
  LAYER via2 ;
   RECT 0 0 129.58 70.11 ;
  LAYER metal3 ;
   RECT 0 0 129.58 70.11 ;
  LAYER via3 ;
   RECT 0 0 129.58 70.11 ;
  LAYER metal4 ;
   RECT 0 0 129.58 70.11 ;
 END
END block_341x369_74

MACRO block_126x648_46
 CLASS BLOCK ;
 FOREIGN block_126x648_46 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 47.88 BY 123.12 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 38.095 2.375 38.665 2.945 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 38.095 85.595 38.665 86.165 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 38.095 91.295 38.665 91.865 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 38.095 96.995 38.665 97.565 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 38.095 102.885 38.665 103.455 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 38.095 108.585 38.665 109.155 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 38.095 114.285 38.665 114.855 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 38.095 119.985 38.665 120.555 ;
  END
 END o7
 PIN o8
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 38.095 8.075 38.665 8.645 ;
  END
 END o8
 PIN o9
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 38.095 13.775 38.665 14.345 ;
  END
 END o9
 PIN o10
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 38.095 19.475 38.665 20.045 ;
  END
 END o10
 PIN o11
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 38.095 25.365 38.665 25.935 ;
  END
 END o11
 PIN o12
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 38.095 31.065 38.665 31.635 ;
  END
 END o12
 PIN o13
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 38.095 36.765 38.665 37.335 ;
  END
 END o13
 PIN o14
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 38.095 42.465 38.665 43.035 ;
  END
 END o14
 PIN o15
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 38.095 74.005 38.665 74.575 ;
  END
 END o15
 PIN o16
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 38.095 79.895 38.665 80.465 ;
  END
 END o16
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 1.235 65.075 1.805 65.645 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 1.235 66.405 1.805 66.975 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 7.315 66.215 7.885 66.785 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 1.235 56.905 1.805 57.475 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 38.095 65.455 38.665 66.025 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 1.235 49.495 1.805 50.065 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 1.235 59.565 1.805 60.135 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 1.235 58.235 1.805 58.805 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 38.095 58.425 38.665 58.995 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 38.855 51.775 39.425 52.345 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 38.095 54.815 38.665 55.385 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 1.995 56.525 2.565 57.095 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 1.235 2.755 1.805 3.325 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 1.235 85.215 1.805 85.785 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 1.235 90.915 1.805 91.485 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 1.235 96.615 1.805 97.185 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 1.235 102.315 1.805 102.885 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 1.235 108.205 1.805 108.775 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 1.235 113.905 1.805 114.475 ;
  END
 END i18
 PIN i19
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 1.235 119.605 1.805 120.175 ;
  END
 END i19
 PIN i20
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 1.235 8.455 1.805 9.025 ;
  END
 END i20
 PIN i21
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 1.235 14.155 1.805 14.725 ;
  END
 END i21
 PIN i22
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 1.235 20.045 1.805 20.615 ;
  END
 END i22
 PIN i23
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 1.235 25.745 1.805 26.315 ;
  END
 END i23
 PIN i24
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 1.235 31.445 1.805 32.015 ;
  END
 END i24
 PIN i25
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 1.235 37.145 1.805 37.715 ;
  END
 END i25
 PIN i26
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 1.235 43.035 1.805 43.605 ;
  END
 END i26
 PIN i27
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 1.235 73.625 1.805 74.195 ;
  END
 END i27
 PIN i28
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 1.235 79.325 1.805 79.895 ;
  END
 END i28
 OBS
  LAYER metal1 ;
   RECT 0 0 47.88 123.12 ;
  LAYER via1 ;
   RECT 0 0 47.88 123.12 ;
  LAYER metal2 ;
   RECT 0 0 47.88 123.12 ;
  LAYER via2 ;
   RECT 0 0 47.88 123.12 ;
  LAYER metal3 ;
   RECT 0 0 47.88 123.12 ;
  LAYER via3 ;
   RECT 0 0 47.88 123.12 ;
  LAYER metal4 ;
   RECT 0 0 47.88 123.12 ;
 END
END block_126x648_46

MACRO block_535x945_130
 CLASS BLOCK ;
 FOREIGN block_535x945_130 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 203.3 BY 179.55 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 25.555 3.705 26.125 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 40.945 56.525 41.515 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 50.445 56.525 51.015 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 135.945 56.525 136.515 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 145.445 56.525 146.015 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 154.945 56.525 155.515 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 59.945 56.525 60.515 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 69.445 56.525 70.015 ;
  END
 END o7
 PIN o8
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 78.945 56.525 79.515 ;
  END
 END o8
 PIN o9
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 88.445 56.525 89.015 ;
  END
 END o9
 PIN o10
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 97.945 56.525 98.515 ;
  END
 END o10
 PIN o11
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 107.445 56.525 108.015 ;
  END
 END o11
 PIN o12
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 116.945 56.525 117.515 ;
  END
 END o12
 PIN o13
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 126.445 56.525 127.015 ;
  END
 END o13
 PIN o14
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 37.715 56.525 38.285 ;
  END
 END o14
 PIN o15
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 47.215 56.525 47.785 ;
  END
 END o15
 PIN o16
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 132.715 56.525 133.285 ;
  END
 END o16
 PIN o17
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 142.215 56.525 142.785 ;
  END
 END o17
 PIN o18
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 151.715 56.525 152.285 ;
  END
 END o18
 PIN o19
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 56.715 56.525 57.285 ;
  END
 END o19
 PIN o20
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 66.215 56.525 66.785 ;
  END
 END o20
 PIN o21
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 75.715 56.525 76.285 ;
  END
 END o21
 PIN o22
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 85.215 56.525 85.785 ;
  END
 END o22
 PIN o23
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 94.715 56.525 95.285 ;
  END
 END o23
 PIN o24
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 104.215 56.525 104.785 ;
  END
 END o24
 PIN o25
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 113.715 56.525 114.285 ;
  END
 END o25
 PIN o26
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 123.215 56.525 123.785 ;
  END
 END o26
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 18.145 3.705 18.715 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 19.095 3.705 19.665 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 13.395 3.705 13.965 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 16.435 3.705 17.005 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 23.275 3.705 23.845 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 16.055 4.465 16.625 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 5.605 3.705 6.175 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 6.555 3.705 7.125 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 4.655 3.705 5.225 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 44.555 56.525 45.125 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 130.055 56.525 130.625 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 111.055 56.525 111.625 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 54.055 56.525 54.625 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 63.555 56.525 64.125 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 139.555 56.525 140.125 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 120.555 56.525 121.125 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 101.555 56.525 102.125 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 73.055 56.525 73.625 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 82.555 56.525 83.125 ;
  END
 END i18
 PIN i19
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 92.055 56.525 92.625 ;
  END
 END i19
 PIN i20
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 35.055 56.525 35.625 ;
  END
 END i20
 PIN i21
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 149.055 56.525 149.625 ;
  END
 END i21
 PIN i22
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 0.855 3.705 1.425 ;
  END
 END i22
 PIN i23
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 26.125 4.465 26.695 ;
  END
 END i23
 PIN i24
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 156.465 56.525 157.035 ;
  END
 END i24
 PIN i25
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 56.715 156.845 57.285 157.415 ;
  END
 END i25
 PIN i26
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 158.555 56.525 159.125 ;
  END
 END i26
 PIN i27
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 157.225 56.525 157.795 ;
  END
 END i27
 PIN i28
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 56.715 157.795 57.285 158.365 ;
  END
 END i28
 PIN i29
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 30.495 3.705 31.065 ;
  END
 END i29
 PIN i30
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 28.975 3.705 29.545 ;
  END
 END i30
 PIN i31
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 2.375 3.705 2.945 ;
  END
 END i31
 PIN i32
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 1.805 4.465 2.375 ;
  END
 END i32
 PIN i33
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 29.925 4.465 30.495 ;
  END
 END i33
 PIN i34
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 28.025 3.705 28.595 ;
  END
 END i34
 PIN i35
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 2.755 4.465 3.325 ;
  END
 END i35
 PIN i36
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 4.275 4.465 4.845 ;
  END
 END i36
 PIN i37
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 3.705 3.705 4.275 ;
  END
 END i37
 PIN i38
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 4.655 29.545 5.225 30.115 ;
  END
 END i38
 PIN i39
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 13.775 4.465 14.345 ;
  END
 END i39
 PIN i40
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 18.525 4.465 19.095 ;
  END
 END i40
 PIN i41
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 17.575 4.465 18.145 ;
  END
 END i41
 PIN i42
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 23.655 4.465 24.225 ;
  END
 END i42
 PIN i43
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 24.225 3.705 24.795 ;
  END
 END i43
 PIN i44
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 5.225 4.465 5.795 ;
  END
 END i44
 PIN i45
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 6.175 4.465 6.745 ;
  END
 END i45
 PIN i46
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 7.125 4.465 7.695 ;
  END
 END i46
 PIN i47
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 10.925 3.705 11.495 ;
  END
 END i47
 PIN i48
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 26.505 3.705 27.075 ;
  END
 END i48
 PIN i49
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 4.655 1.425 5.225 1.995 ;
  END
 END i49
 PIN i50
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 33.725 56.525 34.295 ;
  END
 END i50
 PIN i51
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 43.225 56.525 43.795 ;
  END
 END i51
 PIN i52
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 128.725 56.525 129.295 ;
  END
 END i52
 PIN i53
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 138.225 56.525 138.795 ;
  END
 END i53
 PIN i54
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 147.725 56.525 148.295 ;
  END
 END i54
 PIN i55
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 52.725 56.525 53.295 ;
  END
 END i55
 PIN i56
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 62.225 56.525 62.795 ;
  END
 END i56
 PIN i57
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 71.725 56.525 72.295 ;
  END
 END i57
 PIN i58
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 81.225 56.525 81.795 ;
  END
 END i58
 PIN i59
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 90.725 56.525 91.295 ;
  END
 END i59
 PIN i60
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 100.225 56.525 100.795 ;
  END
 END i60
 PIN i61
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 109.725 56.525 110.295 ;
  END
 END i61
 PIN i62
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 119.225 56.525 119.795 ;
  END
 END i62
 PIN i63
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 38.855 56.525 39.425 ;
  END
 END i63
 PIN i64
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 48.355 56.525 48.925 ;
  END
 END i64
 PIN i65
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 133.855 56.525 134.425 ;
  END
 END i65
 PIN i66
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 143.355 56.525 143.925 ;
  END
 END i66
 PIN i67
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 152.855 56.525 153.425 ;
  END
 END i67
 PIN i68
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 57.855 56.525 58.425 ;
  END
 END i68
 PIN i69
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 67.355 56.525 67.925 ;
  END
 END i69
 PIN i70
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 76.855 56.525 77.425 ;
  END
 END i70
 PIN i71
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 86.355 56.525 86.925 ;
  END
 END i71
 PIN i72
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 95.855 56.525 96.425 ;
  END
 END i72
 PIN i73
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 105.355 56.525 105.925 ;
  END
 END i73
 PIN i74
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 114.855 56.525 115.425 ;
  END
 END i74
 PIN i75
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 124.355 56.525 124.925 ;
  END
 END i75
 PIN i76
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 56.715 158.935 57.285 159.505 ;
  END
 END i76
 PIN i77
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 39.805 56.525 40.375 ;
  END
 END i77
 PIN i78
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 49.305 56.525 49.875 ;
  END
 END i78
 PIN i79
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 134.805 56.525 135.375 ;
  END
 END i79
 PIN i80
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 144.305 56.525 144.875 ;
  END
 END i80
 PIN i81
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 153.805 56.525 154.375 ;
  END
 END i81
 PIN i82
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 58.805 56.525 59.375 ;
  END
 END i82
 PIN i83
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 68.305 56.525 68.875 ;
  END
 END i83
 PIN i84
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 77.805 56.525 78.375 ;
  END
 END i84
 PIN i85
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 87.305 56.525 87.875 ;
  END
 END i85
 PIN i86
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 96.805 56.525 97.375 ;
  END
 END i86
 PIN i87
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 106.305 56.525 106.875 ;
  END
 END i87
 PIN i88
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 115.805 56.525 116.375 ;
  END
 END i88
 PIN i89
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 125.305 56.525 125.875 ;
  END
 END i89
 PIN i90
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 56.715 34.105 57.285 34.675 ;
  END
 END i90
 PIN i91
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 56.715 43.605 57.285 44.175 ;
  END
 END i91
 PIN i92
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 56.715 129.105 57.285 129.675 ;
  END
 END i92
 PIN i93
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 56.715 138.605 57.285 139.175 ;
  END
 END i93
 PIN i94
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 56.715 148.105 57.285 148.675 ;
  END
 END i94
 PIN i95
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 56.715 53.105 57.285 53.675 ;
  END
 END i95
 PIN i96
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 56.715 62.605 57.285 63.175 ;
  END
 END i96
 PIN i97
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 56.715 72.105 57.285 72.675 ;
  END
 END i97
 PIN i98
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 56.715 81.605 57.285 82.175 ;
  END
 END i98
 PIN i99
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 56.715 91.105 57.285 91.675 ;
  END
 END i99
 PIN i100
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 56.715 100.605 57.285 101.175 ;
  END
 END i100
 PIN i101
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 56.715 110.105 57.285 110.675 ;
  END
 END i101
 PIN i102
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 56.715 119.605 57.285 120.175 ;
  END
 END i102
 OBS
  LAYER metal1 ;
   RECT 0.0 0.0 203.3 1.71 ;
   RECT 0.0 1.71 203.3 3.42 ;
   RECT 0.0 3.42 203.3 5.13 ;
   RECT 0.0 5.13 203.3 6.84 ;
   RECT 0.0 6.84 203.3 8.55 ;
   RECT 0.0 8.55 203.3 10.26 ;
   RECT 0.0 10.26 203.3 11.97 ;
   RECT 0.0 11.97 203.3 13.68 ;
   RECT 0.0 13.68 203.3 15.39 ;
   RECT 0.0 15.39 203.3 17.1 ;
   RECT 0.0 17.1 203.3 18.81 ;
   RECT 0.0 18.81 203.3 20.52 ;
   RECT 0.0 20.52 203.3 22.23 ;
   RECT 0.0 22.23 203.3 23.94 ;
   RECT 0.0 23.94 203.3 25.65 ;
   RECT 0.0 25.65 203.3 27.36 ;
   RECT 0.0 27.36 203.3 29.07 ;
   RECT 0.0 29.07 203.3 30.78 ;
   RECT 0.0 30.78 203.3 32.49 ;
   RECT 0.0 32.49 203.3 34.2 ;
   RECT 52.82 34.2 203.3 35.91 ;
   RECT 52.82 35.91 203.3 37.62 ;
   RECT 52.82 37.62 203.3 39.33 ;
   RECT 52.82 39.33 203.3 41.04 ;
   RECT 52.82 41.04 203.3 42.75 ;
   RECT 52.82 42.75 203.3 44.46 ;
   RECT 52.82 44.46 203.3 46.17 ;
   RECT 52.82 46.17 203.3 47.88 ;
   RECT 52.82 47.88 203.3 49.59 ;
   RECT 52.82 49.59 203.3 51.3 ;
   RECT 52.82 51.3 203.3 53.01 ;
   RECT 52.82 53.01 203.3 54.72 ;
   RECT 52.82 54.72 203.3 56.43 ;
   RECT 52.82 56.43 203.3 58.14 ;
   RECT 52.82 58.14 203.3 59.85 ;
   RECT 52.82 59.85 203.3 61.56 ;
   RECT 52.82 61.56 203.3 63.27 ;
   RECT 52.82 63.27 203.3 64.98 ;
   RECT 52.82 64.98 203.3 66.69 ;
   RECT 52.82 66.69 203.3 68.4 ;
   RECT 52.82 68.4 203.3 70.11 ;
   RECT 52.82 70.11 203.3 71.82 ;
   RECT 52.82 71.82 203.3 73.53 ;
   RECT 52.82 73.53 203.3 75.24 ;
   RECT 52.82 75.24 203.3 76.95 ;
   RECT 52.82 76.95 203.3 78.66 ;
   RECT 52.82 78.66 203.3 80.37 ;
   RECT 52.82 80.37 203.3 82.08 ;
   RECT 52.82 82.08 203.3 83.79 ;
   RECT 52.82 83.79 203.3 85.5 ;
   RECT 52.82 85.5 203.3 87.21 ;
   RECT 52.82 87.21 203.3 88.92 ;
   RECT 52.82 88.92 203.3 90.63 ;
   RECT 52.82 90.63 203.3 92.34 ;
   RECT 52.82 92.34 203.3 94.05 ;
   RECT 52.82 94.05 203.3 95.76 ;
   RECT 52.82 95.76 203.3 97.47 ;
   RECT 52.82 97.47 203.3 99.18 ;
   RECT 52.82 99.18 203.3 100.89 ;
   RECT 52.82 100.89 203.3 102.6 ;
   RECT 52.82 102.6 203.3 104.31 ;
   RECT 52.82 104.31 203.3 106.02 ;
   RECT 52.82 106.02 203.3 107.73 ;
   RECT 52.82 107.73 203.3 109.44 ;
   RECT 52.82 109.44 203.3 111.15 ;
   RECT 52.82 111.15 203.3 112.86 ;
   RECT 52.82 112.86 203.3 114.57 ;
   RECT 52.82 114.57 203.3 116.28 ;
   RECT 52.82 116.28 203.3 117.99 ;
   RECT 52.82 117.99 203.3 119.7 ;
   RECT 52.82 119.7 203.3 121.41 ;
   RECT 52.82 121.41 203.3 123.12 ;
   RECT 52.82 123.12 203.3 124.83 ;
   RECT 52.82 124.83 203.3 126.54 ;
   RECT 52.82 126.54 203.3 128.25 ;
   RECT 52.82 128.25 203.3 129.96 ;
   RECT 52.82 129.96 203.3 131.67 ;
   RECT 52.82 131.67 203.3 133.38 ;
   RECT 52.82 133.38 203.3 135.09 ;
   RECT 52.82 135.09 203.3 136.8 ;
   RECT 52.82 136.8 203.3 138.51 ;
   RECT 52.82 138.51 203.3 140.22 ;
   RECT 52.82 140.22 203.3 141.93 ;
   RECT 52.82 141.93 203.3 143.64 ;
   RECT 52.82 143.64 203.3 145.35 ;
   RECT 52.82 145.35 203.3 147.06 ;
   RECT 52.82 147.06 203.3 148.77 ;
   RECT 52.82 148.77 203.3 150.48 ;
   RECT 52.82 150.48 203.3 152.19 ;
   RECT 52.82 152.19 203.3 153.9 ;
   RECT 52.82 153.9 203.3 155.61 ;
   RECT 52.82 155.61 203.3 157.32 ;
   RECT 52.82 157.32 203.3 159.03 ;
   RECT 52.82 159.03 203.3 160.74 ;
   RECT 52.82 160.74 203.3 162.45 ;
   RECT 52.82 162.45 203.3 164.16 ;
   RECT 52.82 164.16 203.3 165.87 ;
   RECT 52.82 165.87 203.3 167.58 ;
   RECT 52.82 167.58 203.3 169.29 ;
   RECT 52.82 169.29 203.3 171.0 ;
   RECT 52.82 171.0 203.3 172.71 ;
   RECT 52.82 172.71 203.3 174.42 ;
   RECT 52.82 174.42 203.3 176.13 ;
   RECT 52.82 176.13 203.3 177.84 ;
   RECT 52.82 177.84 203.3 179.55 ;
  LAYER via1 ;
   RECT 0.0 0.0 203.3 1.71 ;
   RECT 0.0 1.71 203.3 3.42 ;
   RECT 0.0 3.42 203.3 5.13 ;
   RECT 0.0 5.13 203.3 6.84 ;
   RECT 0.0 6.84 203.3 8.55 ;
   RECT 0.0 8.55 203.3 10.26 ;
   RECT 0.0 10.26 203.3 11.97 ;
   RECT 0.0 11.97 203.3 13.68 ;
   RECT 0.0 13.68 203.3 15.39 ;
   RECT 0.0 15.39 203.3 17.1 ;
   RECT 0.0 17.1 203.3 18.81 ;
   RECT 0.0 18.81 203.3 20.52 ;
   RECT 0.0 20.52 203.3 22.23 ;
   RECT 0.0 22.23 203.3 23.94 ;
   RECT 0.0 23.94 203.3 25.65 ;
   RECT 0.0 25.65 203.3 27.36 ;
   RECT 0.0 27.36 203.3 29.07 ;
   RECT 0.0 29.07 203.3 30.78 ;
   RECT 0.0 30.78 203.3 32.49 ;
   RECT 0.0 32.49 203.3 34.2 ;
   RECT 52.82 34.2 203.3 35.91 ;
   RECT 52.82 35.91 203.3 37.62 ;
   RECT 52.82 37.62 203.3 39.33 ;
   RECT 52.82 39.33 203.3 41.04 ;
   RECT 52.82 41.04 203.3 42.75 ;
   RECT 52.82 42.75 203.3 44.46 ;
   RECT 52.82 44.46 203.3 46.17 ;
   RECT 52.82 46.17 203.3 47.88 ;
   RECT 52.82 47.88 203.3 49.59 ;
   RECT 52.82 49.59 203.3 51.3 ;
   RECT 52.82 51.3 203.3 53.01 ;
   RECT 52.82 53.01 203.3 54.72 ;
   RECT 52.82 54.72 203.3 56.43 ;
   RECT 52.82 56.43 203.3 58.14 ;
   RECT 52.82 58.14 203.3 59.85 ;
   RECT 52.82 59.85 203.3 61.56 ;
   RECT 52.82 61.56 203.3 63.27 ;
   RECT 52.82 63.27 203.3 64.98 ;
   RECT 52.82 64.98 203.3 66.69 ;
   RECT 52.82 66.69 203.3 68.4 ;
   RECT 52.82 68.4 203.3 70.11 ;
   RECT 52.82 70.11 203.3 71.82 ;
   RECT 52.82 71.82 203.3 73.53 ;
   RECT 52.82 73.53 203.3 75.24 ;
   RECT 52.82 75.24 203.3 76.95 ;
   RECT 52.82 76.95 203.3 78.66 ;
   RECT 52.82 78.66 203.3 80.37 ;
   RECT 52.82 80.37 203.3 82.08 ;
   RECT 52.82 82.08 203.3 83.79 ;
   RECT 52.82 83.79 203.3 85.5 ;
   RECT 52.82 85.5 203.3 87.21 ;
   RECT 52.82 87.21 203.3 88.92 ;
   RECT 52.82 88.92 203.3 90.63 ;
   RECT 52.82 90.63 203.3 92.34 ;
   RECT 52.82 92.34 203.3 94.05 ;
   RECT 52.82 94.05 203.3 95.76 ;
   RECT 52.82 95.76 203.3 97.47 ;
   RECT 52.82 97.47 203.3 99.18 ;
   RECT 52.82 99.18 203.3 100.89 ;
   RECT 52.82 100.89 203.3 102.6 ;
   RECT 52.82 102.6 203.3 104.31 ;
   RECT 52.82 104.31 203.3 106.02 ;
   RECT 52.82 106.02 203.3 107.73 ;
   RECT 52.82 107.73 203.3 109.44 ;
   RECT 52.82 109.44 203.3 111.15 ;
   RECT 52.82 111.15 203.3 112.86 ;
   RECT 52.82 112.86 203.3 114.57 ;
   RECT 52.82 114.57 203.3 116.28 ;
   RECT 52.82 116.28 203.3 117.99 ;
   RECT 52.82 117.99 203.3 119.7 ;
   RECT 52.82 119.7 203.3 121.41 ;
   RECT 52.82 121.41 203.3 123.12 ;
   RECT 52.82 123.12 203.3 124.83 ;
   RECT 52.82 124.83 203.3 126.54 ;
   RECT 52.82 126.54 203.3 128.25 ;
   RECT 52.82 128.25 203.3 129.96 ;
   RECT 52.82 129.96 203.3 131.67 ;
   RECT 52.82 131.67 203.3 133.38 ;
   RECT 52.82 133.38 203.3 135.09 ;
   RECT 52.82 135.09 203.3 136.8 ;
   RECT 52.82 136.8 203.3 138.51 ;
   RECT 52.82 138.51 203.3 140.22 ;
   RECT 52.82 140.22 203.3 141.93 ;
   RECT 52.82 141.93 203.3 143.64 ;
   RECT 52.82 143.64 203.3 145.35 ;
   RECT 52.82 145.35 203.3 147.06 ;
   RECT 52.82 147.06 203.3 148.77 ;
   RECT 52.82 148.77 203.3 150.48 ;
   RECT 52.82 150.48 203.3 152.19 ;
   RECT 52.82 152.19 203.3 153.9 ;
   RECT 52.82 153.9 203.3 155.61 ;
   RECT 52.82 155.61 203.3 157.32 ;
   RECT 52.82 157.32 203.3 159.03 ;
   RECT 52.82 159.03 203.3 160.74 ;
   RECT 52.82 160.74 203.3 162.45 ;
   RECT 52.82 162.45 203.3 164.16 ;
   RECT 52.82 164.16 203.3 165.87 ;
   RECT 52.82 165.87 203.3 167.58 ;
   RECT 52.82 167.58 203.3 169.29 ;
   RECT 52.82 169.29 203.3 171.0 ;
   RECT 52.82 171.0 203.3 172.71 ;
   RECT 52.82 172.71 203.3 174.42 ;
   RECT 52.82 174.42 203.3 176.13 ;
   RECT 52.82 176.13 203.3 177.84 ;
   RECT 52.82 177.84 203.3 179.55 ;
  LAYER metal2 ;
   RECT 0.0 0.0 203.3 1.71 ;
   RECT 0.0 1.71 203.3 3.42 ;
   RECT 0.0 3.42 203.3 5.13 ;
   RECT 0.0 5.13 203.3 6.84 ;
   RECT 0.0 6.84 203.3 8.55 ;
   RECT 0.0 8.55 203.3 10.26 ;
   RECT 0.0 10.26 203.3 11.97 ;
   RECT 0.0 11.97 203.3 13.68 ;
   RECT 0.0 13.68 203.3 15.39 ;
   RECT 0.0 15.39 203.3 17.1 ;
   RECT 0.0 17.1 203.3 18.81 ;
   RECT 0.0 18.81 203.3 20.52 ;
   RECT 0.0 20.52 203.3 22.23 ;
   RECT 0.0 22.23 203.3 23.94 ;
   RECT 0.0 23.94 203.3 25.65 ;
   RECT 0.0 25.65 203.3 27.36 ;
   RECT 0.0 27.36 203.3 29.07 ;
   RECT 0.0 29.07 203.3 30.78 ;
   RECT 0.0 30.78 203.3 32.49 ;
   RECT 0.0 32.49 203.3 34.2 ;
   RECT 52.82 34.2 203.3 35.91 ;
   RECT 52.82 35.91 203.3 37.62 ;
   RECT 52.82 37.62 203.3 39.33 ;
   RECT 52.82 39.33 203.3 41.04 ;
   RECT 52.82 41.04 203.3 42.75 ;
   RECT 52.82 42.75 203.3 44.46 ;
   RECT 52.82 44.46 203.3 46.17 ;
   RECT 52.82 46.17 203.3 47.88 ;
   RECT 52.82 47.88 203.3 49.59 ;
   RECT 52.82 49.59 203.3 51.3 ;
   RECT 52.82 51.3 203.3 53.01 ;
   RECT 52.82 53.01 203.3 54.72 ;
   RECT 52.82 54.72 203.3 56.43 ;
   RECT 52.82 56.43 203.3 58.14 ;
   RECT 52.82 58.14 203.3 59.85 ;
   RECT 52.82 59.85 203.3 61.56 ;
   RECT 52.82 61.56 203.3 63.27 ;
   RECT 52.82 63.27 203.3 64.98 ;
   RECT 52.82 64.98 203.3 66.69 ;
   RECT 52.82 66.69 203.3 68.4 ;
   RECT 52.82 68.4 203.3 70.11 ;
   RECT 52.82 70.11 203.3 71.82 ;
   RECT 52.82 71.82 203.3 73.53 ;
   RECT 52.82 73.53 203.3 75.24 ;
   RECT 52.82 75.24 203.3 76.95 ;
   RECT 52.82 76.95 203.3 78.66 ;
   RECT 52.82 78.66 203.3 80.37 ;
   RECT 52.82 80.37 203.3 82.08 ;
   RECT 52.82 82.08 203.3 83.79 ;
   RECT 52.82 83.79 203.3 85.5 ;
   RECT 52.82 85.5 203.3 87.21 ;
   RECT 52.82 87.21 203.3 88.92 ;
   RECT 52.82 88.92 203.3 90.63 ;
   RECT 52.82 90.63 203.3 92.34 ;
   RECT 52.82 92.34 203.3 94.05 ;
   RECT 52.82 94.05 203.3 95.76 ;
   RECT 52.82 95.76 203.3 97.47 ;
   RECT 52.82 97.47 203.3 99.18 ;
   RECT 52.82 99.18 203.3 100.89 ;
   RECT 52.82 100.89 203.3 102.6 ;
   RECT 52.82 102.6 203.3 104.31 ;
   RECT 52.82 104.31 203.3 106.02 ;
   RECT 52.82 106.02 203.3 107.73 ;
   RECT 52.82 107.73 203.3 109.44 ;
   RECT 52.82 109.44 203.3 111.15 ;
   RECT 52.82 111.15 203.3 112.86 ;
   RECT 52.82 112.86 203.3 114.57 ;
   RECT 52.82 114.57 203.3 116.28 ;
   RECT 52.82 116.28 203.3 117.99 ;
   RECT 52.82 117.99 203.3 119.7 ;
   RECT 52.82 119.7 203.3 121.41 ;
   RECT 52.82 121.41 203.3 123.12 ;
   RECT 52.82 123.12 203.3 124.83 ;
   RECT 52.82 124.83 203.3 126.54 ;
   RECT 52.82 126.54 203.3 128.25 ;
   RECT 52.82 128.25 203.3 129.96 ;
   RECT 52.82 129.96 203.3 131.67 ;
   RECT 52.82 131.67 203.3 133.38 ;
   RECT 52.82 133.38 203.3 135.09 ;
   RECT 52.82 135.09 203.3 136.8 ;
   RECT 52.82 136.8 203.3 138.51 ;
   RECT 52.82 138.51 203.3 140.22 ;
   RECT 52.82 140.22 203.3 141.93 ;
   RECT 52.82 141.93 203.3 143.64 ;
   RECT 52.82 143.64 203.3 145.35 ;
   RECT 52.82 145.35 203.3 147.06 ;
   RECT 52.82 147.06 203.3 148.77 ;
   RECT 52.82 148.77 203.3 150.48 ;
   RECT 52.82 150.48 203.3 152.19 ;
   RECT 52.82 152.19 203.3 153.9 ;
   RECT 52.82 153.9 203.3 155.61 ;
   RECT 52.82 155.61 203.3 157.32 ;
   RECT 52.82 157.32 203.3 159.03 ;
   RECT 52.82 159.03 203.3 160.74 ;
   RECT 52.82 160.74 203.3 162.45 ;
   RECT 52.82 162.45 203.3 164.16 ;
   RECT 52.82 164.16 203.3 165.87 ;
   RECT 52.82 165.87 203.3 167.58 ;
   RECT 52.82 167.58 203.3 169.29 ;
   RECT 52.82 169.29 203.3 171.0 ;
   RECT 52.82 171.0 203.3 172.71 ;
   RECT 52.82 172.71 203.3 174.42 ;
   RECT 52.82 174.42 203.3 176.13 ;
   RECT 52.82 176.13 203.3 177.84 ;
   RECT 52.82 177.84 203.3 179.55 ;
  LAYER via2 ;
   RECT 0.0 0.0 203.3 1.71 ;
   RECT 0.0 1.71 203.3 3.42 ;
   RECT 0.0 3.42 203.3 5.13 ;
   RECT 0.0 5.13 203.3 6.84 ;
   RECT 0.0 6.84 203.3 8.55 ;
   RECT 0.0 8.55 203.3 10.26 ;
   RECT 0.0 10.26 203.3 11.97 ;
   RECT 0.0 11.97 203.3 13.68 ;
   RECT 0.0 13.68 203.3 15.39 ;
   RECT 0.0 15.39 203.3 17.1 ;
   RECT 0.0 17.1 203.3 18.81 ;
   RECT 0.0 18.81 203.3 20.52 ;
   RECT 0.0 20.52 203.3 22.23 ;
   RECT 0.0 22.23 203.3 23.94 ;
   RECT 0.0 23.94 203.3 25.65 ;
   RECT 0.0 25.65 203.3 27.36 ;
   RECT 0.0 27.36 203.3 29.07 ;
   RECT 0.0 29.07 203.3 30.78 ;
   RECT 0.0 30.78 203.3 32.49 ;
   RECT 0.0 32.49 203.3 34.2 ;
   RECT 52.82 34.2 203.3 35.91 ;
   RECT 52.82 35.91 203.3 37.62 ;
   RECT 52.82 37.62 203.3 39.33 ;
   RECT 52.82 39.33 203.3 41.04 ;
   RECT 52.82 41.04 203.3 42.75 ;
   RECT 52.82 42.75 203.3 44.46 ;
   RECT 52.82 44.46 203.3 46.17 ;
   RECT 52.82 46.17 203.3 47.88 ;
   RECT 52.82 47.88 203.3 49.59 ;
   RECT 52.82 49.59 203.3 51.3 ;
   RECT 52.82 51.3 203.3 53.01 ;
   RECT 52.82 53.01 203.3 54.72 ;
   RECT 52.82 54.72 203.3 56.43 ;
   RECT 52.82 56.43 203.3 58.14 ;
   RECT 52.82 58.14 203.3 59.85 ;
   RECT 52.82 59.85 203.3 61.56 ;
   RECT 52.82 61.56 203.3 63.27 ;
   RECT 52.82 63.27 203.3 64.98 ;
   RECT 52.82 64.98 203.3 66.69 ;
   RECT 52.82 66.69 203.3 68.4 ;
   RECT 52.82 68.4 203.3 70.11 ;
   RECT 52.82 70.11 203.3 71.82 ;
   RECT 52.82 71.82 203.3 73.53 ;
   RECT 52.82 73.53 203.3 75.24 ;
   RECT 52.82 75.24 203.3 76.95 ;
   RECT 52.82 76.95 203.3 78.66 ;
   RECT 52.82 78.66 203.3 80.37 ;
   RECT 52.82 80.37 203.3 82.08 ;
   RECT 52.82 82.08 203.3 83.79 ;
   RECT 52.82 83.79 203.3 85.5 ;
   RECT 52.82 85.5 203.3 87.21 ;
   RECT 52.82 87.21 203.3 88.92 ;
   RECT 52.82 88.92 203.3 90.63 ;
   RECT 52.82 90.63 203.3 92.34 ;
   RECT 52.82 92.34 203.3 94.05 ;
   RECT 52.82 94.05 203.3 95.76 ;
   RECT 52.82 95.76 203.3 97.47 ;
   RECT 52.82 97.47 203.3 99.18 ;
   RECT 52.82 99.18 203.3 100.89 ;
   RECT 52.82 100.89 203.3 102.6 ;
   RECT 52.82 102.6 203.3 104.31 ;
   RECT 52.82 104.31 203.3 106.02 ;
   RECT 52.82 106.02 203.3 107.73 ;
   RECT 52.82 107.73 203.3 109.44 ;
   RECT 52.82 109.44 203.3 111.15 ;
   RECT 52.82 111.15 203.3 112.86 ;
   RECT 52.82 112.86 203.3 114.57 ;
   RECT 52.82 114.57 203.3 116.28 ;
   RECT 52.82 116.28 203.3 117.99 ;
   RECT 52.82 117.99 203.3 119.7 ;
   RECT 52.82 119.7 203.3 121.41 ;
   RECT 52.82 121.41 203.3 123.12 ;
   RECT 52.82 123.12 203.3 124.83 ;
   RECT 52.82 124.83 203.3 126.54 ;
   RECT 52.82 126.54 203.3 128.25 ;
   RECT 52.82 128.25 203.3 129.96 ;
   RECT 52.82 129.96 203.3 131.67 ;
   RECT 52.82 131.67 203.3 133.38 ;
   RECT 52.82 133.38 203.3 135.09 ;
   RECT 52.82 135.09 203.3 136.8 ;
   RECT 52.82 136.8 203.3 138.51 ;
   RECT 52.82 138.51 203.3 140.22 ;
   RECT 52.82 140.22 203.3 141.93 ;
   RECT 52.82 141.93 203.3 143.64 ;
   RECT 52.82 143.64 203.3 145.35 ;
   RECT 52.82 145.35 203.3 147.06 ;
   RECT 52.82 147.06 203.3 148.77 ;
   RECT 52.82 148.77 203.3 150.48 ;
   RECT 52.82 150.48 203.3 152.19 ;
   RECT 52.82 152.19 203.3 153.9 ;
   RECT 52.82 153.9 203.3 155.61 ;
   RECT 52.82 155.61 203.3 157.32 ;
   RECT 52.82 157.32 203.3 159.03 ;
   RECT 52.82 159.03 203.3 160.74 ;
   RECT 52.82 160.74 203.3 162.45 ;
   RECT 52.82 162.45 203.3 164.16 ;
   RECT 52.82 164.16 203.3 165.87 ;
   RECT 52.82 165.87 203.3 167.58 ;
   RECT 52.82 167.58 203.3 169.29 ;
   RECT 52.82 169.29 203.3 171.0 ;
   RECT 52.82 171.0 203.3 172.71 ;
   RECT 52.82 172.71 203.3 174.42 ;
   RECT 52.82 174.42 203.3 176.13 ;
   RECT 52.82 176.13 203.3 177.84 ;
   RECT 52.82 177.84 203.3 179.55 ;
  LAYER metal3 ;
   RECT 0.0 0.0 203.3 1.71 ;
   RECT 0.0 1.71 203.3 3.42 ;
   RECT 0.0 3.42 203.3 5.13 ;
   RECT 0.0 5.13 203.3 6.84 ;
   RECT 0.0 6.84 203.3 8.55 ;
   RECT 0.0 8.55 203.3 10.26 ;
   RECT 0.0 10.26 203.3 11.97 ;
   RECT 0.0 11.97 203.3 13.68 ;
   RECT 0.0 13.68 203.3 15.39 ;
   RECT 0.0 15.39 203.3 17.1 ;
   RECT 0.0 17.1 203.3 18.81 ;
   RECT 0.0 18.81 203.3 20.52 ;
   RECT 0.0 20.52 203.3 22.23 ;
   RECT 0.0 22.23 203.3 23.94 ;
   RECT 0.0 23.94 203.3 25.65 ;
   RECT 0.0 25.65 203.3 27.36 ;
   RECT 0.0 27.36 203.3 29.07 ;
   RECT 0.0 29.07 203.3 30.78 ;
   RECT 0.0 30.78 203.3 32.49 ;
   RECT 0.0 32.49 203.3 34.2 ;
   RECT 52.82 34.2 203.3 35.91 ;
   RECT 52.82 35.91 203.3 37.62 ;
   RECT 52.82 37.62 203.3 39.33 ;
   RECT 52.82 39.33 203.3 41.04 ;
   RECT 52.82 41.04 203.3 42.75 ;
   RECT 52.82 42.75 203.3 44.46 ;
   RECT 52.82 44.46 203.3 46.17 ;
   RECT 52.82 46.17 203.3 47.88 ;
   RECT 52.82 47.88 203.3 49.59 ;
   RECT 52.82 49.59 203.3 51.3 ;
   RECT 52.82 51.3 203.3 53.01 ;
   RECT 52.82 53.01 203.3 54.72 ;
   RECT 52.82 54.72 203.3 56.43 ;
   RECT 52.82 56.43 203.3 58.14 ;
   RECT 52.82 58.14 203.3 59.85 ;
   RECT 52.82 59.85 203.3 61.56 ;
   RECT 52.82 61.56 203.3 63.27 ;
   RECT 52.82 63.27 203.3 64.98 ;
   RECT 52.82 64.98 203.3 66.69 ;
   RECT 52.82 66.69 203.3 68.4 ;
   RECT 52.82 68.4 203.3 70.11 ;
   RECT 52.82 70.11 203.3 71.82 ;
   RECT 52.82 71.82 203.3 73.53 ;
   RECT 52.82 73.53 203.3 75.24 ;
   RECT 52.82 75.24 203.3 76.95 ;
   RECT 52.82 76.95 203.3 78.66 ;
   RECT 52.82 78.66 203.3 80.37 ;
   RECT 52.82 80.37 203.3 82.08 ;
   RECT 52.82 82.08 203.3 83.79 ;
   RECT 52.82 83.79 203.3 85.5 ;
   RECT 52.82 85.5 203.3 87.21 ;
   RECT 52.82 87.21 203.3 88.92 ;
   RECT 52.82 88.92 203.3 90.63 ;
   RECT 52.82 90.63 203.3 92.34 ;
   RECT 52.82 92.34 203.3 94.05 ;
   RECT 52.82 94.05 203.3 95.76 ;
   RECT 52.82 95.76 203.3 97.47 ;
   RECT 52.82 97.47 203.3 99.18 ;
   RECT 52.82 99.18 203.3 100.89 ;
   RECT 52.82 100.89 203.3 102.6 ;
   RECT 52.82 102.6 203.3 104.31 ;
   RECT 52.82 104.31 203.3 106.02 ;
   RECT 52.82 106.02 203.3 107.73 ;
   RECT 52.82 107.73 203.3 109.44 ;
   RECT 52.82 109.44 203.3 111.15 ;
   RECT 52.82 111.15 203.3 112.86 ;
   RECT 52.82 112.86 203.3 114.57 ;
   RECT 52.82 114.57 203.3 116.28 ;
   RECT 52.82 116.28 203.3 117.99 ;
   RECT 52.82 117.99 203.3 119.7 ;
   RECT 52.82 119.7 203.3 121.41 ;
   RECT 52.82 121.41 203.3 123.12 ;
   RECT 52.82 123.12 203.3 124.83 ;
   RECT 52.82 124.83 203.3 126.54 ;
   RECT 52.82 126.54 203.3 128.25 ;
   RECT 52.82 128.25 203.3 129.96 ;
   RECT 52.82 129.96 203.3 131.67 ;
   RECT 52.82 131.67 203.3 133.38 ;
   RECT 52.82 133.38 203.3 135.09 ;
   RECT 52.82 135.09 203.3 136.8 ;
   RECT 52.82 136.8 203.3 138.51 ;
   RECT 52.82 138.51 203.3 140.22 ;
   RECT 52.82 140.22 203.3 141.93 ;
   RECT 52.82 141.93 203.3 143.64 ;
   RECT 52.82 143.64 203.3 145.35 ;
   RECT 52.82 145.35 203.3 147.06 ;
   RECT 52.82 147.06 203.3 148.77 ;
   RECT 52.82 148.77 203.3 150.48 ;
   RECT 52.82 150.48 203.3 152.19 ;
   RECT 52.82 152.19 203.3 153.9 ;
   RECT 52.82 153.9 203.3 155.61 ;
   RECT 52.82 155.61 203.3 157.32 ;
   RECT 52.82 157.32 203.3 159.03 ;
   RECT 52.82 159.03 203.3 160.74 ;
   RECT 52.82 160.74 203.3 162.45 ;
   RECT 52.82 162.45 203.3 164.16 ;
   RECT 52.82 164.16 203.3 165.87 ;
   RECT 52.82 165.87 203.3 167.58 ;
   RECT 52.82 167.58 203.3 169.29 ;
   RECT 52.82 169.29 203.3 171.0 ;
   RECT 52.82 171.0 203.3 172.71 ;
   RECT 52.82 172.71 203.3 174.42 ;
   RECT 52.82 174.42 203.3 176.13 ;
   RECT 52.82 176.13 203.3 177.84 ;
   RECT 52.82 177.84 203.3 179.55 ;
  LAYER via3 ;
   RECT 0.0 0.0 203.3 1.71 ;
   RECT 0.0 1.71 203.3 3.42 ;
   RECT 0.0 3.42 203.3 5.13 ;
   RECT 0.0 5.13 203.3 6.84 ;
   RECT 0.0 6.84 203.3 8.55 ;
   RECT 0.0 8.55 203.3 10.26 ;
   RECT 0.0 10.26 203.3 11.97 ;
   RECT 0.0 11.97 203.3 13.68 ;
   RECT 0.0 13.68 203.3 15.39 ;
   RECT 0.0 15.39 203.3 17.1 ;
   RECT 0.0 17.1 203.3 18.81 ;
   RECT 0.0 18.81 203.3 20.52 ;
   RECT 0.0 20.52 203.3 22.23 ;
   RECT 0.0 22.23 203.3 23.94 ;
   RECT 0.0 23.94 203.3 25.65 ;
   RECT 0.0 25.65 203.3 27.36 ;
   RECT 0.0 27.36 203.3 29.07 ;
   RECT 0.0 29.07 203.3 30.78 ;
   RECT 0.0 30.78 203.3 32.49 ;
   RECT 0.0 32.49 203.3 34.2 ;
   RECT 52.82 34.2 203.3 35.91 ;
   RECT 52.82 35.91 203.3 37.62 ;
   RECT 52.82 37.62 203.3 39.33 ;
   RECT 52.82 39.33 203.3 41.04 ;
   RECT 52.82 41.04 203.3 42.75 ;
   RECT 52.82 42.75 203.3 44.46 ;
   RECT 52.82 44.46 203.3 46.17 ;
   RECT 52.82 46.17 203.3 47.88 ;
   RECT 52.82 47.88 203.3 49.59 ;
   RECT 52.82 49.59 203.3 51.3 ;
   RECT 52.82 51.3 203.3 53.01 ;
   RECT 52.82 53.01 203.3 54.72 ;
   RECT 52.82 54.72 203.3 56.43 ;
   RECT 52.82 56.43 203.3 58.14 ;
   RECT 52.82 58.14 203.3 59.85 ;
   RECT 52.82 59.85 203.3 61.56 ;
   RECT 52.82 61.56 203.3 63.27 ;
   RECT 52.82 63.27 203.3 64.98 ;
   RECT 52.82 64.98 203.3 66.69 ;
   RECT 52.82 66.69 203.3 68.4 ;
   RECT 52.82 68.4 203.3 70.11 ;
   RECT 52.82 70.11 203.3 71.82 ;
   RECT 52.82 71.82 203.3 73.53 ;
   RECT 52.82 73.53 203.3 75.24 ;
   RECT 52.82 75.24 203.3 76.95 ;
   RECT 52.82 76.95 203.3 78.66 ;
   RECT 52.82 78.66 203.3 80.37 ;
   RECT 52.82 80.37 203.3 82.08 ;
   RECT 52.82 82.08 203.3 83.79 ;
   RECT 52.82 83.79 203.3 85.5 ;
   RECT 52.82 85.5 203.3 87.21 ;
   RECT 52.82 87.21 203.3 88.92 ;
   RECT 52.82 88.92 203.3 90.63 ;
   RECT 52.82 90.63 203.3 92.34 ;
   RECT 52.82 92.34 203.3 94.05 ;
   RECT 52.82 94.05 203.3 95.76 ;
   RECT 52.82 95.76 203.3 97.47 ;
   RECT 52.82 97.47 203.3 99.18 ;
   RECT 52.82 99.18 203.3 100.89 ;
   RECT 52.82 100.89 203.3 102.6 ;
   RECT 52.82 102.6 203.3 104.31 ;
   RECT 52.82 104.31 203.3 106.02 ;
   RECT 52.82 106.02 203.3 107.73 ;
   RECT 52.82 107.73 203.3 109.44 ;
   RECT 52.82 109.44 203.3 111.15 ;
   RECT 52.82 111.15 203.3 112.86 ;
   RECT 52.82 112.86 203.3 114.57 ;
   RECT 52.82 114.57 203.3 116.28 ;
   RECT 52.82 116.28 203.3 117.99 ;
   RECT 52.82 117.99 203.3 119.7 ;
   RECT 52.82 119.7 203.3 121.41 ;
   RECT 52.82 121.41 203.3 123.12 ;
   RECT 52.82 123.12 203.3 124.83 ;
   RECT 52.82 124.83 203.3 126.54 ;
   RECT 52.82 126.54 203.3 128.25 ;
   RECT 52.82 128.25 203.3 129.96 ;
   RECT 52.82 129.96 203.3 131.67 ;
   RECT 52.82 131.67 203.3 133.38 ;
   RECT 52.82 133.38 203.3 135.09 ;
   RECT 52.82 135.09 203.3 136.8 ;
   RECT 52.82 136.8 203.3 138.51 ;
   RECT 52.82 138.51 203.3 140.22 ;
   RECT 52.82 140.22 203.3 141.93 ;
   RECT 52.82 141.93 203.3 143.64 ;
   RECT 52.82 143.64 203.3 145.35 ;
   RECT 52.82 145.35 203.3 147.06 ;
   RECT 52.82 147.06 203.3 148.77 ;
   RECT 52.82 148.77 203.3 150.48 ;
   RECT 52.82 150.48 203.3 152.19 ;
   RECT 52.82 152.19 203.3 153.9 ;
   RECT 52.82 153.9 203.3 155.61 ;
   RECT 52.82 155.61 203.3 157.32 ;
   RECT 52.82 157.32 203.3 159.03 ;
   RECT 52.82 159.03 203.3 160.74 ;
   RECT 52.82 160.74 203.3 162.45 ;
   RECT 52.82 162.45 203.3 164.16 ;
   RECT 52.82 164.16 203.3 165.87 ;
   RECT 52.82 165.87 203.3 167.58 ;
   RECT 52.82 167.58 203.3 169.29 ;
   RECT 52.82 169.29 203.3 171.0 ;
   RECT 52.82 171.0 203.3 172.71 ;
   RECT 52.82 172.71 203.3 174.42 ;
   RECT 52.82 174.42 203.3 176.13 ;
   RECT 52.82 176.13 203.3 177.84 ;
   RECT 52.82 177.84 203.3 179.55 ;
  LAYER metal4 ;
   RECT 0.0 0.0 203.3 1.71 ;
   RECT 0.0 1.71 203.3 3.42 ;
   RECT 0.0 3.42 203.3 5.13 ;
   RECT 0.0 5.13 203.3 6.84 ;
   RECT 0.0 6.84 203.3 8.55 ;
   RECT 0.0 8.55 203.3 10.26 ;
   RECT 0.0 10.26 203.3 11.97 ;
   RECT 0.0 11.97 203.3 13.68 ;
   RECT 0.0 13.68 203.3 15.39 ;
   RECT 0.0 15.39 203.3 17.1 ;
   RECT 0.0 17.1 203.3 18.81 ;
   RECT 0.0 18.81 203.3 20.52 ;
   RECT 0.0 20.52 203.3 22.23 ;
   RECT 0.0 22.23 203.3 23.94 ;
   RECT 0.0 23.94 203.3 25.65 ;
   RECT 0.0 25.65 203.3 27.36 ;
   RECT 0.0 27.36 203.3 29.07 ;
   RECT 0.0 29.07 203.3 30.78 ;
   RECT 0.0 30.78 203.3 32.49 ;
   RECT 0.0 32.49 203.3 34.2 ;
   RECT 52.82 34.2 203.3 35.91 ;
   RECT 52.82 35.91 203.3 37.62 ;
   RECT 52.82 37.62 203.3 39.33 ;
   RECT 52.82 39.33 203.3 41.04 ;
   RECT 52.82 41.04 203.3 42.75 ;
   RECT 52.82 42.75 203.3 44.46 ;
   RECT 52.82 44.46 203.3 46.17 ;
   RECT 52.82 46.17 203.3 47.88 ;
   RECT 52.82 47.88 203.3 49.59 ;
   RECT 52.82 49.59 203.3 51.3 ;
   RECT 52.82 51.3 203.3 53.01 ;
   RECT 52.82 53.01 203.3 54.72 ;
   RECT 52.82 54.72 203.3 56.43 ;
   RECT 52.82 56.43 203.3 58.14 ;
   RECT 52.82 58.14 203.3 59.85 ;
   RECT 52.82 59.85 203.3 61.56 ;
   RECT 52.82 61.56 203.3 63.27 ;
   RECT 52.82 63.27 203.3 64.98 ;
   RECT 52.82 64.98 203.3 66.69 ;
   RECT 52.82 66.69 203.3 68.4 ;
   RECT 52.82 68.4 203.3 70.11 ;
   RECT 52.82 70.11 203.3 71.82 ;
   RECT 52.82 71.82 203.3 73.53 ;
   RECT 52.82 73.53 203.3 75.24 ;
   RECT 52.82 75.24 203.3 76.95 ;
   RECT 52.82 76.95 203.3 78.66 ;
   RECT 52.82 78.66 203.3 80.37 ;
   RECT 52.82 80.37 203.3 82.08 ;
   RECT 52.82 82.08 203.3 83.79 ;
   RECT 52.82 83.79 203.3 85.5 ;
   RECT 52.82 85.5 203.3 87.21 ;
   RECT 52.82 87.21 203.3 88.92 ;
   RECT 52.82 88.92 203.3 90.63 ;
   RECT 52.82 90.63 203.3 92.34 ;
   RECT 52.82 92.34 203.3 94.05 ;
   RECT 52.82 94.05 203.3 95.76 ;
   RECT 52.82 95.76 203.3 97.47 ;
   RECT 52.82 97.47 203.3 99.18 ;
   RECT 52.82 99.18 203.3 100.89 ;
   RECT 52.82 100.89 203.3 102.6 ;
   RECT 52.82 102.6 203.3 104.31 ;
   RECT 52.82 104.31 203.3 106.02 ;
   RECT 52.82 106.02 203.3 107.73 ;
   RECT 52.82 107.73 203.3 109.44 ;
   RECT 52.82 109.44 203.3 111.15 ;
   RECT 52.82 111.15 203.3 112.86 ;
   RECT 52.82 112.86 203.3 114.57 ;
   RECT 52.82 114.57 203.3 116.28 ;
   RECT 52.82 116.28 203.3 117.99 ;
   RECT 52.82 117.99 203.3 119.7 ;
   RECT 52.82 119.7 203.3 121.41 ;
   RECT 52.82 121.41 203.3 123.12 ;
   RECT 52.82 123.12 203.3 124.83 ;
   RECT 52.82 124.83 203.3 126.54 ;
   RECT 52.82 126.54 203.3 128.25 ;
   RECT 52.82 128.25 203.3 129.96 ;
   RECT 52.82 129.96 203.3 131.67 ;
   RECT 52.82 131.67 203.3 133.38 ;
   RECT 52.82 133.38 203.3 135.09 ;
   RECT 52.82 135.09 203.3 136.8 ;
   RECT 52.82 136.8 203.3 138.51 ;
   RECT 52.82 138.51 203.3 140.22 ;
   RECT 52.82 140.22 203.3 141.93 ;
   RECT 52.82 141.93 203.3 143.64 ;
   RECT 52.82 143.64 203.3 145.35 ;
   RECT 52.82 145.35 203.3 147.06 ;
   RECT 52.82 147.06 203.3 148.77 ;
   RECT 52.82 148.77 203.3 150.48 ;
   RECT 52.82 150.48 203.3 152.19 ;
   RECT 52.82 152.19 203.3 153.9 ;
   RECT 52.82 153.9 203.3 155.61 ;
   RECT 52.82 155.61 203.3 157.32 ;
   RECT 52.82 157.32 203.3 159.03 ;
   RECT 52.82 159.03 203.3 160.74 ;
   RECT 52.82 160.74 203.3 162.45 ;
   RECT 52.82 162.45 203.3 164.16 ;
   RECT 52.82 164.16 203.3 165.87 ;
   RECT 52.82 165.87 203.3 167.58 ;
   RECT 52.82 167.58 203.3 169.29 ;
   RECT 52.82 169.29 203.3 171.0 ;
   RECT 52.82 171.0 203.3 172.71 ;
   RECT 52.82 172.71 203.3 174.42 ;
   RECT 52.82 174.42 203.3 176.13 ;
   RECT 52.82 176.13 203.3 177.84 ;
   RECT 52.82 177.84 203.3 179.55 ;
 END
END block_535x945_130

MACRO block_546x675_105
 CLASS BLOCK ;
 FOREIGN block_546x675_105 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 207.48 BY 128.25 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 122.835 126.825 123.405 127.395 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 4.275 3.325 4.845 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 20.995 3.325 21.565 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 20.235 3.325 20.805 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 18.715 3.325 19.285 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 62.035 3.325 62.605 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 58.995 3.325 59.565 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 58.235 3.325 58.805 ;
  END
 END o7
 PIN o8
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 18.335 204.345 18.905 ;
  END
 END o8
 PIN o9
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 19.855 204.345 20.425 ;
  END
 END o9
 PIN o10
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 20.615 204.345 21.185 ;
  END
 END o10
 PIN o11
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 21.375 204.345 21.945 ;
  END
 END o11
 PIN o12
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 22.135 204.345 22.705 ;
  END
 END o12
 PIN o13
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 22.895 204.345 23.465 ;
  END
 END o13
 PIN o14
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 24.415 204.345 24.985 ;
  END
 END o14
 PIN o15
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 25.175 204.345 25.745 ;
  END
 END o15
 PIN o16
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 25.935 204.345 26.505 ;
  END
 END o16
 PIN o17
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 26.695 204.345 27.265 ;
  END
 END o17
 PIN o18
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 27.455 204.345 28.025 ;
  END
 END o18
 PIN o19
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 28.975 204.345 29.545 ;
  END
 END o19
 PIN o20
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 29.735 204.345 30.305 ;
  END
 END o20
 PIN o21
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 30.495 204.345 31.065 ;
  END
 END o21
 PIN o22
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 31.255 204.345 31.825 ;
  END
 END o22
 PIN o23
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 48.735 204.345 49.305 ;
  END
 END o23
 PIN o24
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 33.535 204.345 34.105 ;
  END
 END o24
 PIN o25
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 34.295 204.345 34.865 ;
  END
 END o25
 PIN o26
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 35.055 204.345 35.625 ;
  END
 END o26
 PIN o27
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 35.815 204.345 36.385 ;
  END
 END o27
 PIN o28
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 36.575 204.345 37.145 ;
  END
 END o28
 PIN o29
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 38.095 204.345 38.665 ;
  END
 END o29
 PIN o30
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 38.855 204.345 39.425 ;
  END
 END o30
 PIN o31
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 39.615 204.345 40.185 ;
  END
 END o31
 PIN o32
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 40.375 204.345 40.945 ;
  END
 END o32
 PIN o33
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 41.135 204.345 41.705 ;
  END
 END o33
 PIN o34
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 42.655 204.345 43.225 ;
  END
 END o34
 PIN o35
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 43.415 204.345 43.985 ;
  END
 END o35
 PIN o36
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 44.175 204.345 44.745 ;
  END
 END o36
 PIN o37
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 44.935 204.345 45.505 ;
  END
 END o37
 PIN o38
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 45.695 204.345 46.265 ;
  END
 END o38
 PIN o39
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 47.215 204.345 47.785 ;
  END
 END o39
 PIN o40
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 47.975 204.345 48.545 ;
  END
 END o40
 PIN o41
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 49.495 204.345 50.065 ;
  END
 END o41
 PIN o42
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 50.255 204.345 50.825 ;
  END
 END o42
 PIN o43
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 51.775 204.345 52.345 ;
  END
 END o43
 PIN o44
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 52.535 204.345 53.105 ;
  END
 END o44
 PIN o45
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 53.295 204.345 53.865 ;
  END
 END o45
 PIN o46
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 54.055 204.345 54.625 ;
  END
 END o46
 PIN o47
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 54.815 204.345 55.385 ;
  END
 END o47
 PIN o48
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 95.095 126.825 95.665 127.395 ;
  END
 END o48
 PIN o49
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 101.555 126.825 102.125 127.395 ;
  END
 END o49
 PIN o50
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 104.215 126.825 104.785 127.395 ;
  END
 END o50
 PIN o51
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 107.255 126.825 107.825 127.395 ;
  END
 END o51
 PIN o52
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 110.675 126.825 111.245 127.395 ;
  END
 END o52
 PIN o53
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 114.095 126.825 114.665 127.395 ;
  END
 END o53
 PIN o54
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.135 126.825 117.705 127.395 ;
  END
 END o54
 PIN o55
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 119.795 126.825 120.365 127.395 ;
  END
 END o55
 PIN o56
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 132.715 126.825 133.285 127.395 ;
  END
 END o56
 PIN o57
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 153.995 126.825 154.565 127.395 ;
  END
 END o57
 PIN o58
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 172.995 126.825 173.565 127.395 ;
  END
 END o58
 PIN o59
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 176.035 126.825 176.605 127.395 ;
  END
 END o59
 PIN o60
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 179.455 126.825 180.025 127.395 ;
  END
 END o60
 PIN o61
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 181.735 126.825 182.305 127.395 ;
  END
 END o61
 PIN o62
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 185.155 126.825 185.725 127.395 ;
  END
 END o62
 PIN o63
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 188.575 126.825 189.145 127.395 ;
  END
 END o63
 PIN o64
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 191.615 126.825 192.185 127.395 ;
  END
 END o64
 PIN o65
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 200.735 126.825 201.305 127.395 ;
  END
 END o65
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 82.935 126.825 83.505 127.395 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 70.395 126.825 70.965 127.395 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 85.975 126.825 86.545 127.395 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 80.275 3.325 80.845 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 41.895 126.825 42.465 127.395 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 44.935 126.825 45.505 127.395 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 48.355 126.825 48.925 127.395 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 51.775 126.825 52.345 127.395 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 54.815 126.825 55.385 127.395 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 57.475 126.825 58.045 127.395 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 60.515 126.825 61.085 127.395 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 63.935 126.825 64.505 127.395 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 88.635 126.825 89.205 127.395 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 73.055 126.825 73.625 127.395 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 91.675 126.825 92.245 127.395 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 98.515 126.825 99.085 127.395 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 126.825 130.245 127.395 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 150.955 126.825 151.525 127.395 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 197.315 126.825 197.885 127.395 ;
  END
 END i18
 PIN i19
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 56.335 204.345 56.905 ;
  END
 END i19
 PIN i20
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 57.095 204.345 57.665 ;
  END
 END i20
 PIN i21
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 57.855 204.345 58.425 ;
  END
 END i21
 PIN i22
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 58.615 204.345 59.185 ;
  END
 END i22
 PIN i23
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 59.375 204.345 59.945 ;
  END
 END i23
 PIN i24
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 60.895 204.345 61.465 ;
  END
 END i24
 PIN i25
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 61.655 204.345 62.225 ;
  END
 END i25
 PIN i26
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 63.175 204.345 63.745 ;
  END
 END i26
 PIN i27
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 63.935 204.345 64.505 ;
  END
 END i27
 PIN i28
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 65.455 204.345 66.025 ;
  END
 END i28
 PIN i29
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 66.215 204.345 66.785 ;
  END
 END i29
 PIN i30
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 66.975 204.345 67.545 ;
  END
 END i30
 PIN i31
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 67.735 204.345 68.305 ;
  END
 END i31
 PIN i32
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 68.495 204.345 69.065 ;
  END
 END i32
 PIN i33
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 74.955 3.325 75.525 ;
  END
 END i33
 PIN i34
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 75.715 3.325 76.285 ;
  END
 END i34
 PIN i35
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 76.475 3.325 77.045 ;
  END
 END i35
 PIN i36
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 77.235 3.325 77.805 ;
  END
 END i36
 PIN i37
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 77.995 3.325 78.565 ;
  END
 END i37
 PIN i38
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 79.515 3.325 80.085 ;
  END
 END i38
 OBS
  LAYER metal1 ;
   RECT 0 0 207.48 128.25 ;
  LAYER via1 ;
   RECT 0 0 207.48 128.25 ;
  LAYER metal2 ;
   RECT 0 0 207.48 128.25 ;
  LAYER via2 ;
   RECT 0 0 207.48 128.25 ;
  LAYER metal3 ;
   RECT 0 0 207.48 128.25 ;
  LAYER via3 ;
   RECT 0 0 207.48 128.25 ;
  LAYER metal4 ;
   RECT 0 0 207.48 128.25 ;
 END
END block_546x675_105

MACRO block_197x171_33
 CLASS BLOCK ;
 FOREIGN block_197x171_33 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 74.86 BY 32.49 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 25.175 71.725 25.745 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 16.815 71.725 17.385 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 15.295 3.325 15.865 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 16.055 3.325 16.625 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 16.815 3.325 17.385 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 17.575 3.325 18.145 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 18.335 3.325 18.905 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 12.635 3.325 13.205 ;
  END
 END o7
 PIN o8
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 18.335 71.725 18.905 ;
  END
 END o8
 PIN o9
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 9.595 3.325 10.165 ;
  END
 END o9
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 21.375 71.725 21.945 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 70.395 21.755 70.965 22.325 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 22.135 71.725 22.705 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 70.395 22.515 70.965 23.085 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 24.415 71.725 24.985 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 70.395 24.795 70.965 25.365 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 26.695 71.725 27.265 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 27.455 71.725 28.025 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 5.035 3.325 5.605 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 16.055 71.725 16.625 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 13.775 71.725 14.345 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 12.255 71.725 12.825 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 28.975 71.725 29.545 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 25.935 71.725 26.505 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 17.575 71.725 18.145 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 29.735 3.325 30.305 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 22.895 71.725 23.465 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 4.275 71.725 4.845 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 5.035 71.725 5.605 ;
  END
 END i18
 PIN i19
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 6.935 71.725 7.505 ;
  END
 END i19
 PIN i20
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 7.695 71.725 8.265 ;
  END
 END i20
 PIN i21
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 8.835 71.725 9.405 ;
  END
 END i21
 PIN i22
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 9.595 71.725 10.165 ;
  END
 END i22
 OBS
  LAYER metal1 ;
   RECT 0 0 74.86 32.49 ;
  LAYER via1 ;
   RECT 0 0 74.86 32.49 ;
  LAYER metal2 ;
   RECT 0 0 74.86 32.49 ;
  LAYER via2 ;
   RECT 0 0 74.86 32.49 ;
  LAYER metal3 ;
   RECT 0 0 74.86 32.49 ;
  LAYER via3 ;
   RECT 0 0 74.86 32.49 ;
  LAYER metal4 ;
   RECT 0 0 74.86 32.49 ;
 END
END block_197x171_33

MACRO block_2456x4626_834
 CLASS BLOCK ;
 FOREIGN block_2456x4626_834 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 933.28 BY 878.94 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 4.275 26.885 4.845 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 8.455 26.885 9.025 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 45.125 26.885 45.695 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 478.515 26.885 479.085 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 482.695 26.885 483.265 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 486.685 26.885 487.255 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 490.865 26.885 491.435 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 494.855 26.885 495.425 ;
  END
 END o7
 PIN o8
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 499.035 26.885 499.605 ;
  END
 END o8
 PIN o9
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 503.025 26.885 503.595 ;
  END
 END o9
 PIN o10
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 507.205 26.885 507.775 ;
  END
 END o10
 PIN o11
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 511.195 26.885 511.765 ;
  END
 END o11
 PIN o12
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 515.375 26.885 515.945 ;
  END
 END o12
 PIN o13
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 49.305 26.885 49.875 ;
  END
 END o13
 PIN o14
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 519.365 26.885 519.935 ;
  END
 END o14
 PIN o15
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 523.545 26.885 524.115 ;
  END
 END o15
 PIN o16
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 527.535 26.885 528.105 ;
  END
 END o16
 PIN o17
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 531.715 26.885 532.285 ;
  END
 END o17
 PIN o18
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 535.705 26.885 536.275 ;
  END
 END o18
 PIN o19
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 539.885 26.885 540.455 ;
  END
 END o19
 PIN o20
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 543.875 26.885 544.445 ;
  END
 END o20
 PIN o21
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 548.055 26.885 548.625 ;
  END
 END o21
 PIN o22
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 570.285 26.885 570.855 ;
  END
 END o22
 PIN o23
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 574.465 26.885 575.035 ;
  END
 END o23
 PIN o24
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 53.295 26.885 53.865 ;
  END
 END o24
 PIN o25
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 578.455 26.885 579.025 ;
  END
 END o25
 PIN o26
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 582.635 26.885 583.205 ;
  END
 END o26
 PIN o27
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 586.625 26.885 587.195 ;
  END
 END o27
 PIN o28
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 590.805 26.885 591.375 ;
  END
 END o28
 PIN o29
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 594.795 26.885 595.365 ;
  END
 END o29
 PIN o30
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 598.975 26.885 599.545 ;
  END
 END o30
 PIN o31
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 602.965 26.885 603.535 ;
  END
 END o31
 PIN o32
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 607.145 26.885 607.715 ;
  END
 END o32
 PIN o33
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 611.135 26.885 611.705 ;
  END
 END o33
 PIN o34
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 615.315 26.885 615.885 ;
  END
 END o34
 PIN o35
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 57.475 26.885 58.045 ;
  END
 END o35
 PIN o36
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 619.305 26.885 619.875 ;
  END
 END o36
 PIN o37
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 623.485 26.885 624.055 ;
  END
 END o37
 PIN o38
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 627.475 26.885 628.045 ;
  END
 END o38
 PIN o39
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 631.655 26.885 632.225 ;
  END
 END o39
 PIN o40
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 635.645 26.885 636.215 ;
  END
 END o40
 PIN o41
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 639.825 26.885 640.395 ;
  END
 END o41
 PIN o42
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 643.815 26.885 644.385 ;
  END
 END o42
 PIN o43
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 647.995 26.885 648.565 ;
  END
 END o43
 PIN o44
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 651.985 26.885 652.555 ;
  END
 END o44
 PIN o45
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 656.165 26.885 656.735 ;
  END
 END o45
 PIN o46
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 61.465 26.885 62.035 ;
  END
 END o46
 PIN o47
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 660.155 26.885 660.725 ;
  END
 END o47
 PIN o48
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 669.465 26.885 670.035 ;
  END
 END o48
 PIN o49
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 673.455 26.885 674.025 ;
  END
 END o49
 PIN o50
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 677.635 26.885 678.205 ;
  END
 END o50
 PIN o51
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 681.625 26.885 682.195 ;
  END
 END o51
 PIN o52
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 685.805 26.885 686.375 ;
  END
 END o52
 PIN o53
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 689.795 26.885 690.365 ;
  END
 END o53
 PIN o54
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 693.975 26.885 694.545 ;
  END
 END o54
 PIN o55
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 697.965 26.885 698.535 ;
  END
 END o55
 PIN o56
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 702.145 26.885 702.715 ;
  END
 END o56
 PIN o57
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 65.645 26.885 66.215 ;
  END
 END o57
 PIN o58
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 706.135 26.885 706.705 ;
  END
 END o58
 PIN o59
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 710.315 26.885 710.885 ;
  END
 END o59
 PIN o60
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 714.305 26.885 714.875 ;
  END
 END o60
 PIN o61
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 718.485 26.885 719.055 ;
  END
 END o61
 PIN o62
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 722.475 26.885 723.045 ;
  END
 END o62
 PIN o63
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 726.655 26.885 727.225 ;
  END
 END o63
 PIN o64
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 730.645 26.885 731.215 ;
  END
 END o64
 PIN o65
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 734.825 26.885 735.395 ;
  END
 END o65
 PIN o66
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 738.815 26.885 739.385 ;
  END
 END o66
 PIN o67
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 742.995 26.885 743.565 ;
  END
 END o67
 PIN o68
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 69.635 26.885 70.205 ;
  END
 END o68
 PIN o69
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 746.985 26.885 747.555 ;
  END
 END o69
 PIN o70
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 751.165 26.885 751.735 ;
  END
 END o70
 PIN o71
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 755.155 26.885 755.725 ;
  END
 END o71
 PIN o72
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 759.335 26.885 759.905 ;
  END
 END o72
 PIN o73
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 781.565 26.885 782.135 ;
  END
 END o73
 PIN o74
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 785.745 26.885 786.315 ;
  END
 END o74
 PIN o75
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 789.735 26.885 790.305 ;
  END
 END o75
 PIN o76
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 793.915 26.885 794.485 ;
  END
 END o76
 PIN o77
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 797.905 26.885 798.475 ;
  END
 END o77
 PIN o78
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 802.085 26.885 802.655 ;
  END
 END o78
 PIN o79
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 73.815 26.885 74.385 ;
  END
 END o79
 PIN o80
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 806.075 26.885 806.645 ;
  END
 END o80
 PIN o81
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 810.255 26.885 810.825 ;
  END
 END o81
 PIN o82
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 814.245 26.885 814.815 ;
  END
 END o82
 PIN o83
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 818.425 26.885 818.995 ;
  END
 END o83
 PIN o84
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 822.415 26.885 822.985 ;
  END
 END o84
 PIN o85
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 826.595 26.885 827.165 ;
  END
 END o85
 PIN o86
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 830.585 26.885 831.155 ;
  END
 END o86
 PIN o87
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 834.765 26.885 835.335 ;
  END
 END o87
 PIN o88
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 838.755 26.885 839.325 ;
  END
 END o88
 PIN o89
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 842.935 26.885 843.505 ;
  END
 END o89
 PIN o90
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 77.805 26.885 78.375 ;
  END
 END o90
 PIN o91
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 846.925 26.885 847.495 ;
  END
 END o91
 PIN o92
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 851.105 26.885 851.675 ;
  END
 END o92
 PIN o93
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 855.095 26.885 855.665 ;
  END
 END o93
 PIN o94
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 859.275 26.885 859.845 ;
  END
 END o94
 PIN o95
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 863.265 26.885 863.835 ;
  END
 END o95
 PIN o96
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 867.445 26.885 868.015 ;
  END
 END o96
 PIN o97
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 871.435 26.885 872.005 ;
  END
 END o97
 PIN o98
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 81.985 26.885 82.555 ;
  END
 END o98
 PIN o99
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 12.445 26.885 13.015 ;
  END
 END o99
 PIN o100
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 85.975 26.885 86.545 ;
  END
 END o100
 PIN o101
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 90.155 26.885 90.725 ;
  END
 END o101
 PIN o102
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 94.145 26.885 94.715 ;
  END
 END o102
 PIN o103
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 98.325 26.885 98.895 ;
  END
 END o103
 PIN o104
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 120.555 26.885 121.125 ;
  END
 END o104
 PIN o105
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 124.735 26.885 125.305 ;
  END
 END o105
 PIN o106
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 128.725 26.885 129.295 ;
  END
 END o106
 PIN o107
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 132.905 26.885 133.475 ;
  END
 END o107
 PIN o108
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 136.895 26.885 137.465 ;
  END
 END o108
 PIN o109
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 141.075 26.885 141.645 ;
  END
 END o109
 PIN o110
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 16.625 26.885 17.195 ;
  END
 END o110
 PIN o111
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 145.065 26.885 145.635 ;
  END
 END o111
 PIN o112
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 149.245 26.885 149.815 ;
  END
 END o112
 PIN o113
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 153.235 26.885 153.805 ;
  END
 END o113
 PIN o114
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 157.415 26.885 157.985 ;
  END
 END o114
 PIN o115
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 161.405 26.885 161.975 ;
  END
 END o115
 PIN o116
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 165.585 26.885 166.155 ;
  END
 END o116
 PIN o117
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 169.575 26.885 170.145 ;
  END
 END o117
 PIN o118
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 173.755 26.885 174.325 ;
  END
 END o118
 PIN o119
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 177.745 26.885 178.315 ;
  END
 END o119
 PIN o120
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 181.925 26.885 182.495 ;
  END
 END o120
 PIN o121
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 20.615 26.885 21.185 ;
  END
 END o121
 PIN o122
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 185.915 26.885 186.485 ;
  END
 END o122
 PIN o123
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 190.095 26.885 190.665 ;
  END
 END o123
 PIN o124
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 194.085 26.885 194.655 ;
  END
 END o124
 PIN o125
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 198.265 26.885 198.835 ;
  END
 END o125
 PIN o126
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 202.255 26.885 202.825 ;
  END
 END o126
 PIN o127
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 206.435 26.885 207.005 ;
  END
 END o127
 PIN o128
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 210.425 26.885 210.995 ;
  END
 END o128
 PIN o129
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 214.605 26.885 215.175 ;
  END
 END o129
 PIN o130
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 223.725 26.885 224.295 ;
  END
 END o130
 PIN o131
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 227.905 26.885 228.475 ;
  END
 END o131
 PIN o132
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 24.795 26.885 25.365 ;
  END
 END o132
 PIN o133
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 231.895 26.885 232.465 ;
  END
 END o133
 PIN o134
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 236.075 26.885 236.645 ;
  END
 END o134
 PIN o135
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 240.065 26.885 240.635 ;
  END
 END o135
 PIN o136
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 244.245 26.885 244.815 ;
  END
 END o136
 PIN o137
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 248.235 26.885 248.805 ;
  END
 END o137
 PIN o138
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 252.415 26.885 252.985 ;
  END
 END o138
 PIN o139
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 256.405 26.885 256.975 ;
  END
 END o139
 PIN o140
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 260.585 26.885 261.155 ;
  END
 END o140
 PIN o141
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 264.575 26.885 265.145 ;
  END
 END o141
 PIN o142
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 268.755 26.885 269.325 ;
  END
 END o142
 PIN o143
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 28.785 26.885 29.355 ;
  END
 END o143
 PIN o144
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 272.745 26.885 273.315 ;
  END
 END o144
 PIN o145
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 276.925 26.885 277.495 ;
  END
 END o145
 PIN o146
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 280.915 26.885 281.485 ;
  END
 END o146
 PIN o147
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 285.095 26.885 285.665 ;
  END
 END o147
 PIN o148
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 289.085 26.885 289.655 ;
  END
 END o148
 PIN o149
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 293.265 26.885 293.835 ;
  END
 END o149
 PIN o150
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 297.255 26.885 297.825 ;
  END
 END o150
 PIN o151
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 301.435 26.885 302.005 ;
  END
 END o151
 PIN o152
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 305.425 26.885 305.995 ;
  END
 END o152
 PIN o153
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 309.605 26.885 310.175 ;
  END
 END o153
 PIN o154
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 32.965 26.885 33.535 ;
  END
 END o154
 PIN o155
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 313.595 26.885 314.165 ;
  END
 END o155
 PIN o156
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 317.775 26.885 318.345 ;
  END
 END o156
 PIN o157
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 340.005 26.885 340.575 ;
  END
 END o157
 PIN o158
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 344.185 26.885 344.755 ;
  END
 END o158
 PIN o159
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 348.175 26.885 348.745 ;
  END
 END o159
 PIN o160
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 352.355 26.885 352.925 ;
  END
 END o160
 PIN o161
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 356.345 26.885 356.915 ;
  END
 END o161
 PIN o162
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 360.525 26.885 361.095 ;
  END
 END o162
 PIN o163
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 364.515 26.885 365.085 ;
  END
 END o163
 PIN o164
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 368.695 26.885 369.265 ;
  END
 END o164
 PIN o165
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 36.955 26.885 37.525 ;
  END
 END o165
 PIN o166
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 372.685 26.885 373.255 ;
  END
 END o166
 PIN o167
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 376.865 26.885 377.435 ;
  END
 END o167
 PIN o168
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 380.855 26.885 381.425 ;
  END
 END o168
 PIN o169
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 385.035 26.885 385.605 ;
  END
 END o169
 PIN o170
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 389.025 26.885 389.595 ;
  END
 END o170
 PIN o171
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 393.205 26.885 393.775 ;
  END
 END o171
 PIN o172
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 397.195 26.885 397.765 ;
  END
 END o172
 PIN o173
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 401.375 26.885 401.945 ;
  END
 END o173
 PIN o174
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 405.365 26.885 405.935 ;
  END
 END o174
 PIN o175
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 409.545 26.885 410.115 ;
  END
 END o175
 PIN o176
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 41.135 26.885 41.705 ;
  END
 END o176
 PIN o177
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 413.535 26.885 414.105 ;
  END
 END o177
 PIN o178
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 417.715 26.885 418.285 ;
  END
 END o178
 PIN o179
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 421.705 26.885 422.275 ;
  END
 END o179
 PIN o180
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 425.885 26.885 426.455 ;
  END
 END o180
 PIN o181
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 429.875 26.885 430.445 ;
  END
 END o181
 PIN o182
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 458.185 26.885 458.755 ;
  END
 END o182
 PIN o183
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 462.175 26.885 462.745 ;
  END
 END o183
 PIN o184
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 466.355 26.885 466.925 ;
  END
 END o184
 PIN o185
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 470.345 26.885 470.915 ;
  END
 END o185
 PIN o186
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 474.525 26.885 475.095 ;
  END
 END o186
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 432.915 3.705 433.485 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 454.575 3.705 455.145 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 454.195 4.465 454.765 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 450.015 3.705 450.585 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 438.235 3.705 438.805 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 433.295 4.465 433.865 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 432.535 4.465 433.105 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 432.155 3.705 432.725 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 441.845 3.705 442.415 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 454.955 4.465 455.525 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 449.635 4.465 450.205 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 446.405 3.705 446.975 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 449.255 3.705 449.825 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 451.345 3.705 451.915 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 453.815 3.705 454.385 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 455.335 3.705 455.905 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 13.015 431.775 13.585 432.345 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 14.155 431.775 14.725 432.345 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 16.055 431.775 16.625 432.345 ;
  END
 END i18
 PIN i19
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 13.015 445.075 13.585 445.645 ;
  END
 END i19
 PIN i20
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 14.155 445.075 14.725 445.645 ;
  END
 END i20
 PIN i21
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 16.055 445.075 16.625 445.645 ;
  END
 END i21
 PIN i22
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 2.565 26.885 3.135 ;
  END
 END i22
 PIN i23
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 6.745 26.885 7.315 ;
  END
 END i23
 PIN i24
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 43.415 26.885 43.985 ;
  END
 END i24
 PIN i25
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 480.225 26.885 480.795 ;
  END
 END i25
 PIN i26
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 484.405 26.885 484.975 ;
  END
 END i26
 PIN i27
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 488.395 26.885 488.965 ;
  END
 END i27
 PIN i28
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 492.575 26.885 493.145 ;
  END
 END i28
 PIN i29
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 496.565 26.885 497.135 ;
  END
 END i29
 PIN i30
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 500.745 26.885 501.315 ;
  END
 END i30
 PIN i31
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 504.735 26.885 505.305 ;
  END
 END i31
 PIN i32
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 508.915 26.885 509.485 ;
  END
 END i32
 PIN i33
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 512.905 26.885 513.475 ;
  END
 END i33
 PIN i34
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 517.085 26.885 517.655 ;
  END
 END i34
 PIN i35
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 47.595 26.885 48.165 ;
  END
 END i35
 PIN i36
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 521.075 26.885 521.645 ;
  END
 END i36
 PIN i37
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 525.255 26.885 525.825 ;
  END
 END i37
 PIN i38
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 529.245 26.885 529.815 ;
  END
 END i38
 PIN i39
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 533.425 26.885 533.995 ;
  END
 END i39
 PIN i40
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 537.415 26.885 537.985 ;
  END
 END i40
 PIN i41
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 541.595 26.885 542.165 ;
  END
 END i41
 PIN i42
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 545.585 26.885 546.155 ;
  END
 END i42
 PIN i43
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 549.765 26.885 550.335 ;
  END
 END i43
 PIN i44
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 571.995 26.885 572.565 ;
  END
 END i44
 PIN i45
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 576.175 26.885 576.745 ;
  END
 END i45
 PIN i46
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 51.585 26.885 52.155 ;
  END
 END i46
 PIN i47
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 580.165 26.885 580.735 ;
  END
 END i47
 PIN i48
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 584.345 26.885 584.915 ;
  END
 END i48
 PIN i49
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 588.335 26.885 588.905 ;
  END
 END i49
 PIN i50
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 592.515 26.885 593.085 ;
  END
 END i50
 PIN i51
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 596.505 26.885 597.075 ;
  END
 END i51
 PIN i52
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 600.685 26.885 601.255 ;
  END
 END i52
 PIN i53
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 604.675 26.885 605.245 ;
  END
 END i53
 PIN i54
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 608.855 26.885 609.425 ;
  END
 END i54
 PIN i55
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 612.845 26.885 613.415 ;
  END
 END i55
 PIN i56
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 617.025 26.885 617.595 ;
  END
 END i56
 PIN i57
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 55.765 26.885 56.335 ;
  END
 END i57
 PIN i58
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 621.015 26.885 621.585 ;
  END
 END i58
 PIN i59
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 625.195 26.885 625.765 ;
  END
 END i59
 PIN i60
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 629.185 26.885 629.755 ;
  END
 END i60
 PIN i61
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 633.365 26.885 633.935 ;
  END
 END i61
 PIN i62
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 637.355 26.885 637.925 ;
  END
 END i62
 PIN i63
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 641.535 26.885 642.105 ;
  END
 END i63
 PIN i64
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 645.525 26.885 646.095 ;
  END
 END i64
 PIN i65
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 649.705 26.885 650.275 ;
  END
 END i65
 PIN i66
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 653.695 26.885 654.265 ;
  END
 END i66
 PIN i67
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 657.875 26.885 658.445 ;
  END
 END i67
 PIN i68
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 59.755 26.885 60.325 ;
  END
 END i68
 PIN i69
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 661.865 26.885 662.435 ;
  END
 END i69
 PIN i70
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 671.175 26.885 671.745 ;
  END
 END i70
 PIN i71
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 675.165 26.885 675.735 ;
  END
 END i71
 PIN i72
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 679.345 26.885 679.915 ;
  END
 END i72
 PIN i73
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 683.335 26.885 683.905 ;
  END
 END i73
 PIN i74
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 687.515 26.885 688.085 ;
  END
 END i74
 PIN i75
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 691.505 26.885 692.075 ;
  END
 END i75
 PIN i76
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 695.685 26.885 696.255 ;
  END
 END i76
 PIN i77
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 699.675 26.885 700.245 ;
  END
 END i77
 PIN i78
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 703.855 26.885 704.425 ;
  END
 END i78
 PIN i79
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 63.935 26.885 64.505 ;
  END
 END i79
 PIN i80
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 707.845 26.885 708.415 ;
  END
 END i80
 PIN i81
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 712.025 26.885 712.595 ;
  END
 END i81
 PIN i82
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 716.015 26.885 716.585 ;
  END
 END i82
 PIN i83
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 720.195 26.885 720.765 ;
  END
 END i83
 PIN i84
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 724.185 26.885 724.755 ;
  END
 END i84
 PIN i85
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 728.365 26.885 728.935 ;
  END
 END i85
 PIN i86
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 732.355 26.885 732.925 ;
  END
 END i86
 PIN i87
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 736.535 26.885 737.105 ;
  END
 END i87
 PIN i88
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 740.525 26.885 741.095 ;
  END
 END i88
 PIN i89
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 744.705 26.885 745.275 ;
  END
 END i89
 PIN i90
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 67.925 26.885 68.495 ;
  END
 END i90
 PIN i91
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 748.695 26.885 749.265 ;
  END
 END i91
 PIN i92
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 752.875 26.885 753.445 ;
  END
 END i92
 PIN i93
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 756.865 26.885 757.435 ;
  END
 END i93
 PIN i94
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 761.045 26.885 761.615 ;
  END
 END i94
 PIN i95
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 783.275 26.885 783.845 ;
  END
 END i95
 PIN i96
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 787.455 26.885 788.025 ;
  END
 END i96
 PIN i97
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 791.445 26.885 792.015 ;
  END
 END i97
 PIN i98
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 795.625 26.885 796.195 ;
  END
 END i98
 PIN i99
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 799.615 26.885 800.185 ;
  END
 END i99
 PIN i100
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 803.795 26.885 804.365 ;
  END
 END i100
 PIN i101
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 72.105 26.885 72.675 ;
  END
 END i101
 PIN i102
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 807.785 26.885 808.355 ;
  END
 END i102
 PIN i103
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 811.965 26.885 812.535 ;
  END
 END i103
 PIN i104
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 815.955 26.885 816.525 ;
  END
 END i104
 PIN i105
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 820.135 26.885 820.705 ;
  END
 END i105
 PIN i106
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 824.125 26.885 824.695 ;
  END
 END i106
 PIN i107
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 828.305 26.885 828.875 ;
  END
 END i107
 PIN i108
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 832.295 26.885 832.865 ;
  END
 END i108
 PIN i109
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 836.475 26.885 837.045 ;
  END
 END i109
 PIN i110
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 840.465 26.885 841.035 ;
  END
 END i110
 PIN i111
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 844.645 26.885 845.215 ;
  END
 END i111
 PIN i112
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 76.095 26.885 76.665 ;
  END
 END i112
 PIN i113
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 848.635 26.885 849.205 ;
  END
 END i113
 PIN i114
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 852.815 26.885 853.385 ;
  END
 END i114
 PIN i115
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 856.805 26.885 857.375 ;
  END
 END i115
 PIN i116
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 860.985 26.885 861.555 ;
  END
 END i116
 PIN i117
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 864.975 26.885 865.545 ;
  END
 END i117
 PIN i118
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 869.155 26.885 869.725 ;
  END
 END i118
 PIN i119
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 873.145 26.885 873.715 ;
  END
 END i119
 PIN i120
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 80.275 26.885 80.845 ;
  END
 END i120
 PIN i121
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 10.735 26.885 11.305 ;
  END
 END i121
 PIN i122
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 84.265 26.885 84.835 ;
  END
 END i122
 PIN i123
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 88.445 26.885 89.015 ;
  END
 END i123
 PIN i124
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 92.435 26.885 93.005 ;
  END
 END i124
 PIN i125
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 96.615 26.885 97.185 ;
  END
 END i125
 PIN i126
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 118.845 26.885 119.415 ;
  END
 END i126
 PIN i127
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 123.025 26.885 123.595 ;
  END
 END i127
 PIN i128
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 127.015 26.885 127.585 ;
  END
 END i128
 PIN i129
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 131.195 26.885 131.765 ;
  END
 END i129
 PIN i130
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 135.185 26.885 135.755 ;
  END
 END i130
 PIN i131
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 139.365 26.885 139.935 ;
  END
 END i131
 PIN i132
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 14.915 26.885 15.485 ;
  END
 END i132
 PIN i133
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 143.355 26.885 143.925 ;
  END
 END i133
 PIN i134
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 147.535 26.885 148.105 ;
  END
 END i134
 PIN i135
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 151.525 26.885 152.095 ;
  END
 END i135
 PIN i136
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 155.705 26.885 156.275 ;
  END
 END i136
 PIN i137
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 159.695 26.885 160.265 ;
  END
 END i137
 PIN i138
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 163.875 26.885 164.445 ;
  END
 END i138
 PIN i139
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 167.865 26.885 168.435 ;
  END
 END i139
 PIN i140
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 172.045 26.885 172.615 ;
  END
 END i140
 PIN i141
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 176.035 26.885 176.605 ;
  END
 END i141
 PIN i142
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 180.215 26.885 180.785 ;
  END
 END i142
 PIN i143
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 18.905 26.885 19.475 ;
  END
 END i143
 PIN i144
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 184.205 26.885 184.775 ;
  END
 END i144
 PIN i145
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 188.385 26.885 188.955 ;
  END
 END i145
 PIN i146
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 192.375 26.885 192.945 ;
  END
 END i146
 PIN i147
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 196.555 26.885 197.125 ;
  END
 END i147
 PIN i148
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 200.545 26.885 201.115 ;
  END
 END i148
 PIN i149
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 204.725 26.885 205.295 ;
  END
 END i149
 PIN i150
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 208.715 26.885 209.285 ;
  END
 END i150
 PIN i151
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 212.895 26.885 213.465 ;
  END
 END i151
 PIN i152
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 222.015 26.885 222.585 ;
  END
 END i152
 PIN i153
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 226.195 26.885 226.765 ;
  END
 END i153
 PIN i154
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 23.085 26.885 23.655 ;
  END
 END i154
 PIN i155
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 230.185 26.885 230.755 ;
  END
 END i155
 PIN i156
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 234.365 26.885 234.935 ;
  END
 END i156
 PIN i157
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 238.355 26.885 238.925 ;
  END
 END i157
 PIN i158
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 242.535 26.885 243.105 ;
  END
 END i158
 PIN i159
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 246.525 26.885 247.095 ;
  END
 END i159
 PIN i160
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 250.705 26.885 251.275 ;
  END
 END i160
 PIN i161
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 254.695 26.885 255.265 ;
  END
 END i161
 PIN i162
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 258.875 26.885 259.445 ;
  END
 END i162
 PIN i163
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 262.865 26.885 263.435 ;
  END
 END i163
 PIN i164
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 267.045 26.885 267.615 ;
  END
 END i164
 PIN i165
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 27.075 26.885 27.645 ;
  END
 END i165
 PIN i166
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 271.035 26.885 271.605 ;
  END
 END i166
 PIN i167
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 275.215 26.885 275.785 ;
  END
 END i167
 PIN i168
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 279.205 26.885 279.775 ;
  END
 END i168
 PIN i169
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 283.385 26.885 283.955 ;
  END
 END i169
 PIN i170
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 287.375 26.885 287.945 ;
  END
 END i170
 PIN i171
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 291.555 26.885 292.125 ;
  END
 END i171
 PIN i172
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 295.545 26.885 296.115 ;
  END
 END i172
 PIN i173
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 299.725 26.885 300.295 ;
  END
 END i173
 PIN i174
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 303.715 26.885 304.285 ;
  END
 END i174
 PIN i175
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 307.895 26.885 308.465 ;
  END
 END i175
 PIN i176
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 31.255 26.885 31.825 ;
  END
 END i176
 PIN i177
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 311.885 26.885 312.455 ;
  END
 END i177
 PIN i178
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 316.065 26.885 316.635 ;
  END
 END i178
 PIN i179
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 338.295 26.885 338.865 ;
  END
 END i179
 PIN i180
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 342.475 26.885 343.045 ;
  END
 END i180
 PIN i181
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 346.465 26.885 347.035 ;
  END
 END i181
 PIN i182
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 350.645 26.885 351.215 ;
  END
 END i182
 PIN i183
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 354.635 26.885 355.205 ;
  END
 END i183
 PIN i184
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 358.815 26.885 359.385 ;
  END
 END i184
 PIN i185
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 362.805 26.885 363.375 ;
  END
 END i185
 PIN i186
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 366.985 26.885 367.555 ;
  END
 END i186
 PIN i187
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 35.245 26.885 35.815 ;
  END
 END i187
 PIN i188
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 370.975 26.885 371.545 ;
  END
 END i188
 PIN i189
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 375.155 26.885 375.725 ;
  END
 END i189
 PIN i190
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 379.145 26.885 379.715 ;
  END
 END i190
 PIN i191
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 383.325 26.885 383.895 ;
  END
 END i191
 PIN i192
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 387.315 26.885 387.885 ;
  END
 END i192
 PIN i193
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 391.495 26.885 392.065 ;
  END
 END i193
 PIN i194
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 395.485 26.885 396.055 ;
  END
 END i194
 PIN i195
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 399.665 26.885 400.235 ;
  END
 END i195
 PIN i196
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 403.655 26.885 404.225 ;
  END
 END i196
 PIN i197
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 407.835 26.885 408.405 ;
  END
 END i197
 PIN i198
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 39.425 26.885 39.995 ;
  END
 END i198
 PIN i199
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 411.825 26.885 412.395 ;
  END
 END i199
 PIN i200
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 416.005 26.885 416.575 ;
  END
 END i200
 PIN i201
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 419.995 26.885 420.565 ;
  END
 END i201
 PIN i202
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 424.175 26.885 424.745 ;
  END
 END i202
 PIN i203
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 428.165 26.885 428.735 ;
  END
 END i203
 PIN i204
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 459.895 26.885 460.465 ;
  END
 END i204
 PIN i205
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 463.885 26.885 464.455 ;
  END
 END i205
 PIN i206
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 468.065 26.885 468.635 ;
  END
 END i206
 PIN i207
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 472.055 26.885 472.625 ;
  END
 END i207
 PIN i208
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 476.235 26.885 476.805 ;
  END
 END i208
 PIN i209
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 74.385 27.645 74.955 ;
  END
 END i209
 PIN i210
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 78.375 27.645 78.945 ;
  END
 END i210
 PIN i211
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 82.555 27.645 83.125 ;
  END
 END i211
 PIN i212
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 62.035 27.645 62.605 ;
  END
 END i212
 PIN i213
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 66.215 27.645 66.785 ;
  END
 END i213
 PIN i214
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 141.645 27.645 142.215 ;
  END
 END i214
 PIN i215
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 145.635 27.645 146.205 ;
  END
 END i215
 PIN i216
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 149.815 27.645 150.385 ;
  END
 END i216
 PIN i217
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 153.805 27.645 154.375 ;
  END
 END i217
 PIN i218
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 157.985 27.645 158.555 ;
  END
 END i218
 PIN i219
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 293.835 27.645 294.405 ;
  END
 END i219
 PIN i220
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 297.825 27.645 298.395 ;
  END
 END i220
 PIN i221
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 302.005 27.645 302.575 ;
  END
 END i221
 PIN i222
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 281.485 27.645 282.055 ;
  END
 END i222
 PIN i223
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 285.665 27.645 286.235 ;
  END
 END i223
 PIN i224
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 361.095 27.645 361.665 ;
  END
 END i224
 PIN i225
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 365.085 27.645 365.655 ;
  END
 END i225
 PIN i226
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 369.265 27.645 369.835 ;
  END
 END i226
 PIN i227
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 373.255 27.645 373.825 ;
  END
 END i227
 PIN i228
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 377.435 27.645 378.005 ;
  END
 END i228
 PIN i229
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 526.965 27.645 527.535 ;
  END
 END i229
 PIN i230
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 522.975 27.645 523.545 ;
  END
 END i230
 PIN i231
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 518.795 27.645 519.365 ;
  END
 END i231
 PIN i232
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 514.805 27.645 515.375 ;
  END
 END i232
 PIN i233
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 510.625 27.645 511.195 ;
  END
 END i233
 PIN i234
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 594.225 27.645 594.795 ;
  END
 END i234
 PIN i235
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 590.235 27.645 590.805 ;
  END
 END i235
 PIN i236
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 586.055 27.645 586.625 ;
  END
 END i236
 PIN i237
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 606.575 27.645 607.145 ;
  END
 END i237
 PIN i238
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 602.395 27.645 602.965 ;
  END
 END i238
 PIN i239
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 738.245 27.645 738.815 ;
  END
 END i239
 PIN i240
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 734.255 27.645 734.825 ;
  END
 END i240
 PIN i241
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 730.075 27.645 730.645 ;
  END
 END i241
 PIN i242
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 726.085 27.645 726.655 ;
  END
 END i242
 PIN i243
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 721.905 27.645 722.475 ;
  END
 END i243
 PIN i244
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 805.505 27.645 806.075 ;
  END
 END i244
 PIN i245
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 801.515 27.645 802.085 ;
  END
 END i245
 PIN i246
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 797.335 27.645 797.905 ;
  END
 END i246
 PIN i247
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 817.855 27.645 818.425 ;
  END
 END i247
 PIN i248
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 813.675 27.645 814.245 ;
  END
 END i248
 PIN i249
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 70.205 27.645 70.775 ;
  END
 END i249
 PIN i250
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 137.465 27.645 138.035 ;
  END
 END i250
 PIN i251
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 289.655 27.645 290.225 ;
  END
 END i251
 PIN i252
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 356.915 27.645 357.485 ;
  END
 END i252
 PIN i253
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 531.145 27.645 531.715 ;
  END
 END i253
 PIN i254
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 598.405 27.645 598.975 ;
  END
 END i254
 PIN i255
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 742.425 27.645 742.995 ;
  END
 END i255
 PIN i256
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 809.685 27.645 810.255 ;
  END
 END i256
 PIN i257
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 17.955 431.775 18.525 432.345 ;
  END
 END i257
 PIN i258
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 17.955 445.075 18.525 445.645 ;
  END
 END i258
 PIN i259
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 3.135 27.645 3.705 ;
  END
 END i259
 PIN i260
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 7.315 27.645 7.885 ;
  END
 END i260
 PIN i261
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 43.985 27.645 44.555 ;
  END
 END i261
 PIN i262
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 479.655 27.645 480.225 ;
  END
 END i262
 PIN i263
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 483.835 27.645 484.405 ;
  END
 END i263
 PIN i264
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 487.825 27.645 488.395 ;
  END
 END i264
 PIN i265
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 492.005 27.645 492.575 ;
  END
 END i265
 PIN i266
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 495.995 27.645 496.565 ;
  END
 END i266
 PIN i267
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 500.175 27.645 500.745 ;
  END
 END i267
 PIN i268
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 504.165 27.645 504.735 ;
  END
 END i268
 PIN i269
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 508.345 27.645 508.915 ;
  END
 END i269
 PIN i270
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 512.335 27.645 512.905 ;
  END
 END i270
 PIN i271
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 516.515 27.645 517.085 ;
  END
 END i271
 PIN i272
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 48.165 27.645 48.735 ;
  END
 END i272
 PIN i273
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 520.505 27.645 521.075 ;
  END
 END i273
 PIN i274
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 524.685 27.645 525.255 ;
  END
 END i274
 PIN i275
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 528.675 27.645 529.245 ;
  END
 END i275
 PIN i276
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 532.855 27.645 533.425 ;
  END
 END i276
 PIN i277
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 536.845 27.645 537.415 ;
  END
 END i277
 PIN i278
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 541.025 27.645 541.595 ;
  END
 END i278
 PIN i279
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 545.015 27.645 545.585 ;
  END
 END i279
 PIN i280
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 549.195 27.645 549.765 ;
  END
 END i280
 PIN i281
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 571.425 27.645 571.995 ;
  END
 END i281
 PIN i282
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 575.605 27.645 576.175 ;
  END
 END i282
 PIN i283
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 52.155 27.645 52.725 ;
  END
 END i283
 PIN i284
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 579.595 27.645 580.165 ;
  END
 END i284
 PIN i285
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 583.775 27.645 584.345 ;
  END
 END i285
 PIN i286
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 587.765 27.645 588.335 ;
  END
 END i286
 PIN i287
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 591.945 27.645 592.515 ;
  END
 END i287
 PIN i288
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 595.935 27.645 596.505 ;
  END
 END i288
 PIN i289
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 600.115 27.645 600.685 ;
  END
 END i289
 PIN i290
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 604.105 27.645 604.675 ;
  END
 END i290
 PIN i291
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 608.285 27.645 608.855 ;
  END
 END i291
 PIN i292
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 612.275 27.645 612.845 ;
  END
 END i292
 PIN i293
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 616.455 27.645 617.025 ;
  END
 END i293
 PIN i294
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 56.335 27.645 56.905 ;
  END
 END i294
 PIN i295
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 620.445 27.645 621.015 ;
  END
 END i295
 PIN i296
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 624.625 27.645 625.195 ;
  END
 END i296
 PIN i297
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 628.615 27.645 629.185 ;
  END
 END i297
 PIN i298
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 632.795 27.645 633.365 ;
  END
 END i298
 PIN i299
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 636.785 27.645 637.355 ;
  END
 END i299
 PIN i300
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 640.965 27.645 641.535 ;
  END
 END i300
 PIN i301
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 644.955 27.645 645.525 ;
  END
 END i301
 PIN i302
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 649.135 27.645 649.705 ;
  END
 END i302
 PIN i303
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 653.125 27.645 653.695 ;
  END
 END i303
 PIN i304
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 657.305 27.645 657.875 ;
  END
 END i304
 PIN i305
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 60.325 27.645 60.895 ;
  END
 END i305
 PIN i306
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 661.295 27.645 661.865 ;
  END
 END i306
 PIN i307
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 670.605 27.645 671.175 ;
  END
 END i307
 PIN i308
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 674.595 27.645 675.165 ;
  END
 END i308
 PIN i309
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 678.775 27.645 679.345 ;
  END
 END i309
 PIN i310
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 682.765 27.645 683.335 ;
  END
 END i310
 PIN i311
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 686.945 27.645 687.515 ;
  END
 END i311
 PIN i312
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 690.935 27.645 691.505 ;
  END
 END i312
 PIN i313
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 695.115 27.645 695.685 ;
  END
 END i313
 PIN i314
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 699.105 27.645 699.675 ;
  END
 END i314
 PIN i315
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 703.285 27.645 703.855 ;
  END
 END i315
 PIN i316
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 64.505 27.645 65.075 ;
  END
 END i316
 PIN i317
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 707.275 27.645 707.845 ;
  END
 END i317
 PIN i318
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 711.455 27.645 712.025 ;
  END
 END i318
 PIN i319
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 715.445 27.645 716.015 ;
  END
 END i319
 PIN i320
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 719.625 27.645 720.195 ;
  END
 END i320
 PIN i321
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 723.615 27.645 724.185 ;
  END
 END i321
 PIN i322
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 727.795 27.645 728.365 ;
  END
 END i322
 PIN i323
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 731.785 27.645 732.355 ;
  END
 END i323
 PIN i324
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 735.965 27.645 736.535 ;
  END
 END i324
 PIN i325
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 739.955 27.645 740.525 ;
  END
 END i325
 PIN i326
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 744.135 27.645 744.705 ;
  END
 END i326
 PIN i327
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 68.495 27.645 69.065 ;
  END
 END i327
 PIN i328
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 748.125 27.645 748.695 ;
  END
 END i328
 PIN i329
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 752.305 27.645 752.875 ;
  END
 END i329
 PIN i330
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 756.295 27.645 756.865 ;
  END
 END i330
 PIN i331
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 760.475 27.645 761.045 ;
  END
 END i331
 PIN i332
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 782.705 27.645 783.275 ;
  END
 END i332
 PIN i333
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 786.885 27.645 787.455 ;
  END
 END i333
 PIN i334
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 790.875 27.645 791.445 ;
  END
 END i334
 PIN i335
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 795.055 27.645 795.625 ;
  END
 END i335
 PIN i336
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 799.045 27.645 799.615 ;
  END
 END i336
 PIN i337
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 803.225 27.645 803.795 ;
  END
 END i337
 PIN i338
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 72.675 27.645 73.245 ;
  END
 END i338
 PIN i339
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 807.215 27.645 807.785 ;
  END
 END i339
 PIN i340
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 811.395 27.645 811.965 ;
  END
 END i340
 PIN i341
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 815.385 27.645 815.955 ;
  END
 END i341
 PIN i342
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 819.565 27.645 820.135 ;
  END
 END i342
 PIN i343
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 823.555 27.645 824.125 ;
  END
 END i343
 PIN i344
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 827.735 27.645 828.305 ;
  END
 END i344
 PIN i345
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 831.725 27.645 832.295 ;
  END
 END i345
 PIN i346
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 835.905 27.645 836.475 ;
  END
 END i346
 PIN i347
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 839.895 27.645 840.465 ;
  END
 END i347
 PIN i348
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 844.075 27.645 844.645 ;
  END
 END i348
 PIN i349
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 76.665 27.645 77.235 ;
  END
 END i349
 PIN i350
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 848.065 27.645 848.635 ;
  END
 END i350
 PIN i351
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 852.245 27.645 852.815 ;
  END
 END i351
 PIN i352
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 856.235 27.645 856.805 ;
  END
 END i352
 PIN i353
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 860.415 27.645 860.985 ;
  END
 END i353
 PIN i354
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 864.405 27.645 864.975 ;
  END
 END i354
 PIN i355
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 868.585 27.645 869.155 ;
  END
 END i355
 PIN i356
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 872.575 27.645 873.145 ;
  END
 END i356
 PIN i357
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 80.845 27.645 81.415 ;
  END
 END i357
 PIN i358
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 11.305 27.645 11.875 ;
  END
 END i358
 PIN i359
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 84.835 27.645 85.405 ;
  END
 END i359
 PIN i360
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 89.015 27.645 89.585 ;
  END
 END i360
 PIN i361
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 93.005 27.645 93.575 ;
  END
 END i361
 PIN i362
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 97.185 27.645 97.755 ;
  END
 END i362
 PIN i363
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 119.415 27.645 119.985 ;
  END
 END i363
 PIN i364
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 123.595 27.645 124.165 ;
  END
 END i364
 PIN i365
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 127.585 27.645 128.155 ;
  END
 END i365
 PIN i366
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 131.765 27.645 132.335 ;
  END
 END i366
 PIN i367
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 135.755 27.645 136.325 ;
  END
 END i367
 PIN i368
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 139.935 27.645 140.505 ;
  END
 END i368
 PIN i369
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 15.485 27.645 16.055 ;
  END
 END i369
 PIN i370
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 143.925 27.645 144.495 ;
  END
 END i370
 PIN i371
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 148.105 27.645 148.675 ;
  END
 END i371
 PIN i372
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 152.095 27.645 152.665 ;
  END
 END i372
 PIN i373
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 156.275 27.645 156.845 ;
  END
 END i373
 PIN i374
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 160.265 27.645 160.835 ;
  END
 END i374
 PIN i375
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 164.445 27.645 165.015 ;
  END
 END i375
 PIN i376
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 168.435 27.645 169.005 ;
  END
 END i376
 PIN i377
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 172.615 27.645 173.185 ;
  END
 END i377
 PIN i378
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 176.605 27.645 177.175 ;
  END
 END i378
 PIN i379
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 180.785 27.645 181.355 ;
  END
 END i379
 PIN i380
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 19.475 27.645 20.045 ;
  END
 END i380
 PIN i381
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 184.775 27.645 185.345 ;
  END
 END i381
 PIN i382
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 188.955 27.645 189.525 ;
  END
 END i382
 PIN i383
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 192.945 27.645 193.515 ;
  END
 END i383
 PIN i384
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 197.125 27.645 197.695 ;
  END
 END i384
 PIN i385
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 201.115 27.645 201.685 ;
  END
 END i385
 PIN i386
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 205.295 27.645 205.865 ;
  END
 END i386
 PIN i387
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 209.285 27.645 209.855 ;
  END
 END i387
 PIN i388
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 213.465 27.645 214.035 ;
  END
 END i388
 PIN i389
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 222.585 27.645 223.155 ;
  END
 END i389
 PIN i390
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 226.765 27.645 227.335 ;
  END
 END i390
 PIN i391
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 23.655 27.645 24.225 ;
  END
 END i391
 PIN i392
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 230.755 27.645 231.325 ;
  END
 END i392
 PIN i393
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 234.935 27.645 235.505 ;
  END
 END i393
 PIN i394
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 238.925 27.645 239.495 ;
  END
 END i394
 PIN i395
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 243.105 27.645 243.675 ;
  END
 END i395
 PIN i396
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 247.095 27.645 247.665 ;
  END
 END i396
 PIN i397
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 251.275 27.645 251.845 ;
  END
 END i397
 PIN i398
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 255.265 27.645 255.835 ;
  END
 END i398
 PIN i399
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 259.445 27.645 260.015 ;
  END
 END i399
 PIN i400
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 263.435 27.645 264.005 ;
  END
 END i400
 PIN i401
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 267.615 27.645 268.185 ;
  END
 END i401
 PIN i402
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 27.645 27.645 28.215 ;
  END
 END i402
 PIN i403
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 271.605 27.645 272.175 ;
  END
 END i403
 PIN i404
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 275.785 27.645 276.355 ;
  END
 END i404
 PIN i405
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 279.775 27.645 280.345 ;
  END
 END i405
 PIN i406
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 283.955 27.645 284.525 ;
  END
 END i406
 PIN i407
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 287.945 27.645 288.515 ;
  END
 END i407
 PIN i408
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 292.125 27.645 292.695 ;
  END
 END i408
 PIN i409
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 296.115 27.645 296.685 ;
  END
 END i409
 PIN i410
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 300.295 27.645 300.865 ;
  END
 END i410
 PIN i411
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 304.285 27.645 304.855 ;
  END
 END i411
 PIN i412
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 308.465 27.645 309.035 ;
  END
 END i412
 PIN i413
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 31.825 27.645 32.395 ;
  END
 END i413
 PIN i414
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 312.455 27.645 313.025 ;
  END
 END i414
 PIN i415
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 316.635 27.645 317.205 ;
  END
 END i415
 PIN i416
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 338.865 27.645 339.435 ;
  END
 END i416
 PIN i417
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 343.045 27.645 343.615 ;
  END
 END i417
 PIN i418
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 347.035 27.645 347.605 ;
  END
 END i418
 PIN i419
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 351.215 27.645 351.785 ;
  END
 END i419
 PIN i420
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 355.205 27.645 355.775 ;
  END
 END i420
 PIN i421
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 359.385 27.645 359.955 ;
  END
 END i421
 PIN i422
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 363.375 27.645 363.945 ;
  END
 END i422
 PIN i423
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 367.555 27.645 368.125 ;
  END
 END i423
 PIN i424
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 35.815 27.645 36.385 ;
  END
 END i424
 PIN i425
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 371.545 27.645 372.115 ;
  END
 END i425
 PIN i426
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 375.725 27.645 376.295 ;
  END
 END i426
 PIN i427
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 379.715 27.645 380.285 ;
  END
 END i427
 PIN i428
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 383.895 27.645 384.465 ;
  END
 END i428
 PIN i429
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 387.885 27.645 388.455 ;
  END
 END i429
 PIN i430
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 392.065 27.645 392.635 ;
  END
 END i430
 PIN i431
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 396.055 27.645 396.625 ;
  END
 END i431
 PIN i432
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 400.235 27.645 400.805 ;
  END
 END i432
 PIN i433
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 404.225 27.645 404.795 ;
  END
 END i433
 PIN i434
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 408.405 27.645 408.975 ;
  END
 END i434
 PIN i435
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 39.995 27.645 40.565 ;
  END
 END i435
 PIN i436
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 412.395 27.645 412.965 ;
  END
 END i436
 PIN i437
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 416.575 27.645 417.145 ;
  END
 END i437
 PIN i438
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 420.565 27.645 421.135 ;
  END
 END i438
 PIN i439
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 424.745 27.645 425.315 ;
  END
 END i439
 PIN i440
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 428.735 27.645 429.305 ;
  END
 END i440
 PIN i441
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 459.325 27.645 459.895 ;
  END
 END i441
 PIN i442
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 463.315 27.645 463.885 ;
  END
 END i442
 PIN i443
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 467.495 27.645 468.065 ;
  END
 END i443
 PIN i444
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 471.485 27.645 472.055 ;
  END
 END i444
 PIN i445
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 475.665 27.645 476.235 ;
  END
 END i445
 PIN i446
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 439.375 3.705 439.945 ;
  END
 END i446
 PIN i447
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 439.755 4.465 440.325 ;
  END
 END i447
 PIN i448
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 3.705 28.405 4.275 ;
  END
 END i448
 PIN i449
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 7.885 28.405 8.455 ;
  END
 END i449
 PIN i450
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 44.555 28.405 45.125 ;
  END
 END i450
 PIN i451
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 479.085 28.405 479.655 ;
  END
 END i451
 PIN i452
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 483.265 28.405 483.835 ;
  END
 END i452
 PIN i453
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 487.255 28.405 487.825 ;
  END
 END i453
 PIN i454
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 491.435 28.405 492.005 ;
  END
 END i454
 PIN i455
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 495.425 28.405 495.995 ;
  END
 END i455
 PIN i456
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 499.605 28.405 500.175 ;
  END
 END i456
 PIN i457
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 503.595 28.405 504.165 ;
  END
 END i457
 PIN i458
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 507.775 28.405 508.345 ;
  END
 END i458
 PIN i459
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 511.765 28.405 512.335 ;
  END
 END i459
 PIN i460
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 515.945 28.405 516.515 ;
  END
 END i460
 PIN i461
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 48.735 28.405 49.305 ;
  END
 END i461
 PIN i462
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 519.935 28.405 520.505 ;
  END
 END i462
 PIN i463
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 524.115 28.405 524.685 ;
  END
 END i463
 PIN i464
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 528.105 28.405 528.675 ;
  END
 END i464
 PIN i465
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 532.285 28.405 532.855 ;
  END
 END i465
 PIN i466
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 536.275 28.405 536.845 ;
  END
 END i466
 PIN i467
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 540.455 28.405 541.025 ;
  END
 END i467
 PIN i468
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 544.445 28.405 545.015 ;
  END
 END i468
 PIN i469
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 548.625 28.405 549.195 ;
  END
 END i469
 PIN i470
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 570.855 28.405 571.425 ;
  END
 END i470
 PIN i471
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 575.035 28.405 575.605 ;
  END
 END i471
 PIN i472
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 52.725 28.405 53.295 ;
  END
 END i472
 PIN i473
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 579.025 28.405 579.595 ;
  END
 END i473
 PIN i474
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 583.205 28.405 583.775 ;
  END
 END i474
 PIN i475
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 587.195 28.405 587.765 ;
  END
 END i475
 PIN i476
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 591.375 28.405 591.945 ;
  END
 END i476
 PIN i477
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 595.365 28.405 595.935 ;
  END
 END i477
 PIN i478
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 599.545 28.405 600.115 ;
  END
 END i478
 PIN i479
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 603.535 28.405 604.105 ;
  END
 END i479
 PIN i480
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 607.715 28.405 608.285 ;
  END
 END i480
 PIN i481
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 611.705 28.405 612.275 ;
  END
 END i481
 PIN i482
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 615.885 28.405 616.455 ;
  END
 END i482
 PIN i483
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 56.905 28.405 57.475 ;
  END
 END i483
 PIN i484
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 619.875 28.405 620.445 ;
  END
 END i484
 PIN i485
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 624.055 28.405 624.625 ;
  END
 END i485
 PIN i486
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 628.045 28.405 628.615 ;
  END
 END i486
 PIN i487
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 632.225 28.405 632.795 ;
  END
 END i487
 PIN i488
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 636.215 28.405 636.785 ;
  END
 END i488
 PIN i489
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 640.395 28.405 640.965 ;
  END
 END i489
 PIN i490
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 644.385 28.405 644.955 ;
  END
 END i490
 PIN i491
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 648.565 28.405 649.135 ;
  END
 END i491
 PIN i492
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 652.555 28.405 653.125 ;
  END
 END i492
 PIN i493
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 656.735 28.405 657.305 ;
  END
 END i493
 PIN i494
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 60.895 28.405 61.465 ;
  END
 END i494
 PIN i495
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 660.725 28.405 661.295 ;
  END
 END i495
 PIN i496
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 670.035 28.405 670.605 ;
  END
 END i496
 PIN i497
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 674.025 28.405 674.595 ;
  END
 END i497
 PIN i498
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 678.205 28.405 678.775 ;
  END
 END i498
 PIN i499
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 682.195 28.405 682.765 ;
  END
 END i499
 PIN i500
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 686.375 28.405 686.945 ;
  END
 END i500
 PIN i501
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 690.365 28.405 690.935 ;
  END
 END i501
 PIN i502
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 694.545 28.405 695.115 ;
  END
 END i502
 PIN i503
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 698.535 28.405 699.105 ;
  END
 END i503
 PIN i504
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 702.715 28.405 703.285 ;
  END
 END i504
 PIN i505
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 65.075 28.405 65.645 ;
  END
 END i505
 PIN i506
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 706.705 28.405 707.275 ;
  END
 END i506
 PIN i507
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 710.885 28.405 711.455 ;
  END
 END i507
 PIN i508
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 714.875 28.405 715.445 ;
  END
 END i508
 PIN i509
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 719.055 28.405 719.625 ;
  END
 END i509
 PIN i510
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 723.045 28.405 723.615 ;
  END
 END i510
 PIN i511
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 727.225 28.405 727.795 ;
  END
 END i511
 PIN i512
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 731.215 28.405 731.785 ;
  END
 END i512
 PIN i513
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 735.395 28.405 735.965 ;
  END
 END i513
 PIN i514
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 739.385 28.405 739.955 ;
  END
 END i514
 PIN i515
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 743.565 28.405 744.135 ;
  END
 END i515
 PIN i516
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 69.065 28.405 69.635 ;
  END
 END i516
 PIN i517
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 747.555 28.405 748.125 ;
  END
 END i517
 PIN i518
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 751.735 28.405 752.305 ;
  END
 END i518
 PIN i519
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 755.725 28.405 756.295 ;
  END
 END i519
 PIN i520
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 759.905 28.405 760.475 ;
  END
 END i520
 PIN i521
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 782.135 28.405 782.705 ;
  END
 END i521
 PIN i522
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 786.315 28.405 786.885 ;
  END
 END i522
 PIN i523
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 790.305 28.405 790.875 ;
  END
 END i523
 PIN i524
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 794.485 28.405 795.055 ;
  END
 END i524
 PIN i525
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 798.475 28.405 799.045 ;
  END
 END i525
 PIN i526
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 802.655 28.405 803.225 ;
  END
 END i526
 PIN i527
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 73.245 28.405 73.815 ;
  END
 END i527
 PIN i528
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 806.645 28.405 807.215 ;
  END
 END i528
 PIN i529
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 810.825 28.405 811.395 ;
  END
 END i529
 PIN i530
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 814.815 28.405 815.385 ;
  END
 END i530
 PIN i531
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 818.995 28.405 819.565 ;
  END
 END i531
 PIN i532
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 822.985 28.405 823.555 ;
  END
 END i532
 PIN i533
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 827.165 28.405 827.735 ;
  END
 END i533
 PIN i534
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 831.155 28.405 831.725 ;
  END
 END i534
 PIN i535
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 835.335 28.405 835.905 ;
  END
 END i535
 PIN i536
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 839.325 28.405 839.895 ;
  END
 END i536
 PIN i537
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 843.505 28.405 844.075 ;
  END
 END i537
 PIN i538
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 77.235 28.405 77.805 ;
  END
 END i538
 PIN i539
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 847.495 28.405 848.065 ;
  END
 END i539
 PIN i540
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 851.675 28.405 852.245 ;
  END
 END i540
 PIN i541
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 855.665 28.405 856.235 ;
  END
 END i541
 PIN i542
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 859.845 28.405 860.415 ;
  END
 END i542
 PIN i543
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 863.835 28.405 864.405 ;
  END
 END i543
 PIN i544
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 868.015 28.405 868.585 ;
  END
 END i544
 PIN i545
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 872.005 28.405 872.575 ;
  END
 END i545
 PIN i546
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 81.415 28.405 81.985 ;
  END
 END i546
 PIN i547
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 11.875 28.405 12.445 ;
  END
 END i547
 PIN i548
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 85.405 28.405 85.975 ;
  END
 END i548
 PIN i549
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 89.585 28.405 90.155 ;
  END
 END i549
 PIN i550
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 93.575 28.405 94.145 ;
  END
 END i550
 PIN i551
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 97.755 28.405 98.325 ;
  END
 END i551
 PIN i552
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 119.985 28.405 120.555 ;
  END
 END i552
 PIN i553
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 124.165 28.405 124.735 ;
  END
 END i553
 PIN i554
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 128.155 28.405 128.725 ;
  END
 END i554
 PIN i555
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 132.335 28.405 132.905 ;
  END
 END i555
 PIN i556
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 136.325 28.405 136.895 ;
  END
 END i556
 PIN i557
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 140.505 28.405 141.075 ;
  END
 END i557
 PIN i558
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 16.055 28.405 16.625 ;
  END
 END i558
 PIN i559
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 144.495 28.405 145.065 ;
  END
 END i559
 PIN i560
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 148.675 28.405 149.245 ;
  END
 END i560
 PIN i561
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 152.665 28.405 153.235 ;
  END
 END i561
 PIN i562
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 156.845 28.405 157.415 ;
  END
 END i562
 PIN i563
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 160.835 28.405 161.405 ;
  END
 END i563
 PIN i564
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 165.015 28.405 165.585 ;
  END
 END i564
 PIN i565
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 169.005 28.405 169.575 ;
  END
 END i565
 PIN i566
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 173.185 28.405 173.755 ;
  END
 END i566
 PIN i567
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 177.175 28.405 177.745 ;
  END
 END i567
 PIN i568
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 181.355 28.405 181.925 ;
  END
 END i568
 PIN i569
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 20.045 28.405 20.615 ;
  END
 END i569
 PIN i570
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 185.345 28.405 185.915 ;
  END
 END i570
 PIN i571
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 189.525 28.405 190.095 ;
  END
 END i571
 PIN i572
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 193.515 28.405 194.085 ;
  END
 END i572
 PIN i573
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 197.695 28.405 198.265 ;
  END
 END i573
 PIN i574
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 201.685 28.405 202.255 ;
  END
 END i574
 PIN i575
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 205.865 28.405 206.435 ;
  END
 END i575
 PIN i576
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 209.855 28.405 210.425 ;
  END
 END i576
 PIN i577
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 214.035 28.405 214.605 ;
  END
 END i577
 PIN i578
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 223.155 28.405 223.725 ;
  END
 END i578
 PIN i579
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 227.335 28.405 227.905 ;
  END
 END i579
 PIN i580
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 24.225 28.405 24.795 ;
  END
 END i580
 PIN i581
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 231.325 28.405 231.895 ;
  END
 END i581
 PIN i582
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 235.505 28.405 236.075 ;
  END
 END i582
 PIN i583
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 239.495 28.405 240.065 ;
  END
 END i583
 PIN i584
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 243.675 28.405 244.245 ;
  END
 END i584
 PIN i585
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 247.665 28.405 248.235 ;
  END
 END i585
 PIN i586
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 251.845 28.405 252.415 ;
  END
 END i586
 PIN i587
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 255.835 28.405 256.405 ;
  END
 END i587
 PIN i588
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 260.015 28.405 260.585 ;
  END
 END i588
 PIN i589
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 264.005 28.405 264.575 ;
  END
 END i589
 PIN i590
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 268.185 28.405 268.755 ;
  END
 END i590
 PIN i591
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 28.215 28.405 28.785 ;
  END
 END i591
 PIN i592
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 272.175 28.405 272.745 ;
  END
 END i592
 PIN i593
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 276.355 28.405 276.925 ;
  END
 END i593
 PIN i594
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 280.345 28.405 280.915 ;
  END
 END i594
 PIN i595
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 284.525 28.405 285.095 ;
  END
 END i595
 PIN i596
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 288.515 28.405 289.085 ;
  END
 END i596
 PIN i597
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 292.695 28.405 293.265 ;
  END
 END i597
 PIN i598
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 296.685 28.405 297.255 ;
  END
 END i598
 PIN i599
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 300.865 28.405 301.435 ;
  END
 END i599
 PIN i600
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 304.855 28.405 305.425 ;
  END
 END i600
 PIN i601
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 309.035 28.405 309.605 ;
  END
 END i601
 PIN i602
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 32.395 28.405 32.965 ;
  END
 END i602
 PIN i603
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 313.025 28.405 313.595 ;
  END
 END i603
 PIN i604
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 317.205 28.405 317.775 ;
  END
 END i604
 PIN i605
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 339.435 28.405 340.005 ;
  END
 END i605
 PIN i606
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 343.615 28.405 344.185 ;
  END
 END i606
 PIN i607
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 347.605 28.405 348.175 ;
  END
 END i607
 PIN i608
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 351.785 28.405 352.355 ;
  END
 END i608
 PIN i609
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 355.775 28.405 356.345 ;
  END
 END i609
 PIN i610
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 359.955 28.405 360.525 ;
  END
 END i610
 PIN i611
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 363.945 28.405 364.515 ;
  END
 END i611
 PIN i612
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 368.125 28.405 368.695 ;
  END
 END i612
 PIN i613
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 36.385 28.405 36.955 ;
  END
 END i613
 PIN i614
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 372.115 28.405 372.685 ;
  END
 END i614
 PIN i615
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 376.295 28.405 376.865 ;
  END
 END i615
 PIN i616
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 380.285 28.405 380.855 ;
  END
 END i616
 PIN i617
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 384.465 28.405 385.035 ;
  END
 END i617
 PIN i618
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 388.455 28.405 389.025 ;
  END
 END i618
 PIN i619
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 392.635 28.405 393.205 ;
  END
 END i619
 PIN i620
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 396.625 28.405 397.195 ;
  END
 END i620
 PIN i621
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 400.805 28.405 401.375 ;
  END
 END i621
 PIN i622
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 404.795 28.405 405.365 ;
  END
 END i622
 PIN i623
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 408.975 28.405 409.545 ;
  END
 END i623
 PIN i624
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 40.565 28.405 41.135 ;
  END
 END i624
 PIN i625
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 412.965 28.405 413.535 ;
  END
 END i625
 PIN i626
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 417.145 28.405 417.715 ;
  END
 END i626
 PIN i627
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 421.135 28.405 421.705 ;
  END
 END i627
 PIN i628
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 425.315 28.405 425.885 ;
  END
 END i628
 PIN i629
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 429.305 28.405 429.875 ;
  END
 END i629
 PIN i630
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 458.755 28.405 459.325 ;
  END
 END i630
 PIN i631
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 462.745 28.405 463.315 ;
  END
 END i631
 PIN i632
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 466.925 28.405 467.495 ;
  END
 END i632
 PIN i633
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 470.915 28.405 471.485 ;
  END
 END i633
 PIN i634
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 475.095 28.405 475.665 ;
  END
 END i634
 PIN i635
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 4.275 431.775 4.845 432.345 ;
  END
 END i635
 PIN i636
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 5.415 431.775 5.985 432.345 ;
  END
 END i636
 PIN i637
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 6.935 431.775 7.505 432.345 ;
  END
 END i637
 PIN i638
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 8.835 431.775 9.405 432.345 ;
  END
 END i638
 PIN i639
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.975 431.775 10.545 432.345 ;
  END
 END i639
 PIN i640
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 11.875 431.775 12.445 432.345 ;
  END
 END i640
 PIN i641
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 4.275 445.075 4.845 445.645 ;
  END
 END i641
 PIN i642
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 5.415 445.075 5.985 445.645 ;
  END
 END i642
 PIN i643
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 6.935 445.075 7.505 445.645 ;
  END
 END i643
 PIN i644
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 8.835 445.075 9.405 445.645 ;
  END
 END i644
 PIN i645
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.975 445.075 10.545 445.645 ;
  END
 END i645
 PIN i646
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 11.875 445.075 12.445 445.645 ;
  END
 END i646
 OBS
  LAYER metal1 ;
   RECT 23.18 0.0 933.28 1.71 ;
   RECT 23.18 1.71 933.28 3.42 ;
   RECT 23.18 3.42 933.28 5.13 ;
   RECT 23.18 5.13 933.28 6.84 ;
   RECT 23.18 6.84 933.28 8.55 ;
   RECT 23.18 8.55 933.28 10.26 ;
   RECT 23.18 10.26 933.28 11.97 ;
   RECT 23.18 11.97 933.28 13.68 ;
   RECT 23.18 13.68 933.28 15.39 ;
   RECT 23.18 15.39 933.28 17.1 ;
   RECT 23.18 17.1 933.28 18.81 ;
   RECT 23.18 18.81 933.28 20.52 ;
   RECT 23.18 20.52 933.28 22.23 ;
   RECT 23.18 22.23 933.28 23.94 ;
   RECT 23.18 23.94 933.28 25.65 ;
   RECT 23.18 25.65 933.28 27.36 ;
   RECT 23.18 27.36 933.28 29.07 ;
   RECT 23.18 29.07 933.28 30.78 ;
   RECT 23.18 30.78 933.28 32.49 ;
   RECT 23.18 32.49 933.28 34.2 ;
   RECT 23.18 34.2 933.28 35.91 ;
   RECT 23.18 35.91 933.28 37.62 ;
   RECT 23.18 37.62 933.28 39.33 ;
   RECT 23.18 39.33 933.28 41.04 ;
   RECT 23.18 41.04 933.28 42.75 ;
   RECT 23.18 42.75 933.28 44.46 ;
   RECT 23.18 44.46 933.28 46.17 ;
   RECT 23.18 46.17 933.28 47.88 ;
   RECT 23.18 47.88 933.28 49.59 ;
   RECT 23.18 49.59 933.28 51.3 ;
   RECT 23.18 51.3 933.28 53.01 ;
   RECT 23.18 53.01 933.28 54.72 ;
   RECT 23.18 54.72 933.28 56.43 ;
   RECT 23.18 56.43 933.28 58.14 ;
   RECT 23.18 58.14 933.28 59.85 ;
   RECT 23.18 59.85 933.28 61.56 ;
   RECT 23.18 61.56 933.28 63.27 ;
   RECT 23.18 63.27 933.28 64.98 ;
   RECT 23.18 64.98 933.28 66.69 ;
   RECT 23.18 66.69 933.28 68.4 ;
   RECT 23.18 68.4 933.28 70.11 ;
   RECT 23.18 70.11 933.28 71.82 ;
   RECT 23.18 71.82 933.28 73.53 ;
   RECT 23.18 73.53 933.28 75.24 ;
   RECT 23.18 75.24 933.28 76.95 ;
   RECT 23.18 76.95 933.28 78.66 ;
   RECT 23.18 78.66 933.28 80.37 ;
   RECT 23.18 80.37 933.28 82.08 ;
   RECT 23.18 82.08 933.28 83.79 ;
   RECT 23.18 83.79 933.28 85.5 ;
   RECT 23.18 85.5 933.28 87.21 ;
   RECT 23.18 87.21 933.28 88.92 ;
   RECT 23.18 88.92 933.28 90.63 ;
   RECT 23.18 90.63 933.28 92.34 ;
   RECT 23.18 92.34 933.28 94.05 ;
   RECT 23.18 94.05 933.28 95.76 ;
   RECT 23.18 95.76 933.28 97.47 ;
   RECT 23.18 97.47 933.28 99.18 ;
   RECT 23.18 99.18 933.28 100.89 ;
   RECT 23.18 100.89 933.28 102.6 ;
   RECT 23.18 102.6 933.28 104.31 ;
   RECT 23.18 104.31 933.28 106.02 ;
   RECT 23.18 106.02 933.28 107.73 ;
   RECT 23.18 107.73 933.28 109.44 ;
   RECT 23.18 109.44 933.28 111.15 ;
   RECT 23.18 111.15 933.28 112.86 ;
   RECT 23.18 112.86 933.28 114.57 ;
   RECT 23.18 114.57 933.28 116.28 ;
   RECT 23.18 116.28 933.28 117.99 ;
   RECT 23.18 117.99 933.28 119.7 ;
   RECT 23.18 119.7 933.28 121.41 ;
   RECT 23.18 121.41 933.28 123.12 ;
   RECT 23.18 123.12 933.28 124.83 ;
   RECT 23.18 124.83 933.28 126.54 ;
   RECT 23.18 126.54 933.28 128.25 ;
   RECT 23.18 128.25 933.28 129.96 ;
   RECT 23.18 129.96 933.28 131.67 ;
   RECT 23.18 131.67 933.28 133.38 ;
   RECT 23.18 133.38 933.28 135.09 ;
   RECT 23.18 135.09 933.28 136.8 ;
   RECT 23.18 136.8 933.28 138.51 ;
   RECT 23.18 138.51 933.28 140.22 ;
   RECT 23.18 140.22 933.28 141.93 ;
   RECT 23.18 141.93 933.28 143.64 ;
   RECT 23.18 143.64 933.28 145.35 ;
   RECT 23.18 145.35 933.28 147.06 ;
   RECT 23.18 147.06 933.28 148.77 ;
   RECT 23.18 148.77 933.28 150.48 ;
   RECT 23.18 150.48 933.28 152.19 ;
   RECT 23.18 152.19 933.28 153.9 ;
   RECT 23.18 153.9 933.28 155.61 ;
   RECT 23.18 155.61 933.28 157.32 ;
   RECT 23.18 157.32 933.28 159.03 ;
   RECT 23.18 159.03 933.28 160.74 ;
   RECT 23.18 160.74 933.28 162.45 ;
   RECT 23.18 162.45 933.28 164.16 ;
   RECT 23.18 164.16 933.28 165.87 ;
   RECT 23.18 165.87 933.28 167.58 ;
   RECT 23.18 167.58 933.28 169.29 ;
   RECT 23.18 169.29 933.28 171.0 ;
   RECT 23.18 171.0 933.28 172.71 ;
   RECT 23.18 172.71 933.28 174.42 ;
   RECT 23.18 174.42 933.28 176.13 ;
   RECT 23.18 176.13 933.28 177.84 ;
   RECT 23.18 177.84 933.28 179.55 ;
   RECT 23.18 179.55 933.28 181.26 ;
   RECT 23.18 181.26 933.28 182.97 ;
   RECT 23.18 182.97 933.28 184.68 ;
   RECT 23.18 184.68 933.28 186.39 ;
   RECT 23.18 186.39 933.28 188.1 ;
   RECT 23.18 188.1 933.28 189.81 ;
   RECT 23.18 189.81 933.28 191.52 ;
   RECT 23.18 191.52 933.28 193.23 ;
   RECT 23.18 193.23 933.28 194.94 ;
   RECT 23.18 194.94 933.28 196.65 ;
   RECT 23.18 196.65 933.28 198.36 ;
   RECT 23.18 198.36 933.28 200.07 ;
   RECT 23.18 200.07 933.28 201.78 ;
   RECT 23.18 201.78 933.28 203.49 ;
   RECT 23.18 203.49 933.28 205.2 ;
   RECT 23.18 205.2 933.28 206.91 ;
   RECT 23.18 206.91 933.28 208.62 ;
   RECT 23.18 208.62 933.28 210.33 ;
   RECT 23.18 210.33 933.28 212.04 ;
   RECT 23.18 212.04 933.28 213.75 ;
   RECT 23.18 213.75 933.28 215.46 ;
   RECT 23.18 215.46 933.28 217.17 ;
   RECT 23.18 217.17 933.28 218.88 ;
   RECT 23.18 218.88 933.28 220.59 ;
   RECT 23.18 220.59 933.28 222.3 ;
   RECT 23.18 222.3 933.28 224.01 ;
   RECT 23.18 224.01 933.28 225.72 ;
   RECT 23.18 225.72 933.28 227.43 ;
   RECT 23.18 227.43 933.28 229.14 ;
   RECT 23.18 229.14 933.28 230.85 ;
   RECT 23.18 230.85 933.28 232.56 ;
   RECT 23.18 232.56 933.28 234.27 ;
   RECT 23.18 234.27 933.28 235.98 ;
   RECT 23.18 235.98 933.28 237.69 ;
   RECT 23.18 237.69 933.28 239.4 ;
   RECT 23.18 239.4 933.28 241.11 ;
   RECT 23.18 241.11 933.28 242.82 ;
   RECT 23.18 242.82 933.28 244.53 ;
   RECT 23.18 244.53 933.28 246.24 ;
   RECT 23.18 246.24 933.28 247.95 ;
   RECT 23.18 247.95 933.28 249.66 ;
   RECT 23.18 249.66 933.28 251.37 ;
   RECT 23.18 251.37 933.28 253.08 ;
   RECT 23.18 253.08 933.28 254.79 ;
   RECT 23.18 254.79 933.28 256.5 ;
   RECT 23.18 256.5 933.28 258.21 ;
   RECT 23.18 258.21 933.28 259.92 ;
   RECT 23.18 259.92 933.28 261.63 ;
   RECT 23.18 261.63 933.28 263.34 ;
   RECT 23.18 263.34 933.28 265.05 ;
   RECT 23.18 265.05 933.28 266.76 ;
   RECT 23.18 266.76 933.28 268.47 ;
   RECT 23.18 268.47 933.28 270.18 ;
   RECT 23.18 270.18 933.28 271.89 ;
   RECT 23.18 271.89 933.28 273.6 ;
   RECT 23.18 273.6 933.28 275.31 ;
   RECT 23.18 275.31 933.28 277.02 ;
   RECT 23.18 277.02 933.28 278.73 ;
   RECT 23.18 278.73 933.28 280.44 ;
   RECT 23.18 280.44 933.28 282.15 ;
   RECT 23.18 282.15 933.28 283.86 ;
   RECT 23.18 283.86 933.28 285.57 ;
   RECT 23.18 285.57 933.28 287.28 ;
   RECT 23.18 287.28 933.28 288.99 ;
   RECT 23.18 288.99 933.28 290.7 ;
   RECT 23.18 290.7 933.28 292.41 ;
   RECT 23.18 292.41 933.28 294.12 ;
   RECT 23.18 294.12 933.28 295.83 ;
   RECT 23.18 295.83 933.28 297.54 ;
   RECT 23.18 297.54 933.28 299.25 ;
   RECT 23.18 299.25 933.28 300.96 ;
   RECT 23.18 300.96 933.28 302.67 ;
   RECT 23.18 302.67 933.28 304.38 ;
   RECT 23.18 304.38 933.28 306.09 ;
   RECT 23.18 306.09 933.28 307.8 ;
   RECT 23.18 307.8 933.28 309.51 ;
   RECT 23.18 309.51 933.28 311.22 ;
   RECT 23.18 311.22 933.28 312.93 ;
   RECT 23.18 312.93 933.28 314.64 ;
   RECT 23.18 314.64 933.28 316.35 ;
   RECT 23.18 316.35 933.28 318.06 ;
   RECT 23.18 318.06 933.28 319.77 ;
   RECT 23.18 319.77 933.28 321.48 ;
   RECT 23.18 321.48 933.28 323.19 ;
   RECT 23.18 323.19 933.28 324.9 ;
   RECT 23.18 324.9 933.28 326.61 ;
   RECT 23.18 326.61 933.28 328.32 ;
   RECT 23.18 328.32 933.28 330.03 ;
   RECT 23.18 330.03 933.28 331.74 ;
   RECT 23.18 331.74 933.28 333.45 ;
   RECT 23.18 333.45 933.28 335.16 ;
   RECT 23.18 335.16 933.28 336.87 ;
   RECT 23.18 336.87 933.28 338.58 ;
   RECT 23.18 338.58 933.28 340.29 ;
   RECT 23.18 340.29 933.28 342.0 ;
   RECT 23.18 342.0 933.28 343.71 ;
   RECT 23.18 343.71 933.28 345.42 ;
   RECT 23.18 345.42 933.28 347.13 ;
   RECT 23.18 347.13 933.28 348.84 ;
   RECT 23.18 348.84 933.28 350.55 ;
   RECT 23.18 350.55 933.28 352.26 ;
   RECT 23.18 352.26 933.28 353.97 ;
   RECT 23.18 353.97 933.28 355.68 ;
   RECT 23.18 355.68 933.28 357.39 ;
   RECT 23.18 357.39 933.28 359.1 ;
   RECT 23.18 359.1 933.28 360.81 ;
   RECT 23.18 360.81 933.28 362.52 ;
   RECT 23.18 362.52 933.28 364.23 ;
   RECT 23.18 364.23 933.28 365.94 ;
   RECT 23.18 365.94 933.28 367.65 ;
   RECT 23.18 367.65 933.28 369.36 ;
   RECT 23.18 369.36 933.28 371.07 ;
   RECT 23.18 371.07 933.28 372.78 ;
   RECT 23.18 372.78 933.28 374.49 ;
   RECT 23.18 374.49 933.28 376.2 ;
   RECT 23.18 376.2 933.28 377.91 ;
   RECT 23.18 377.91 933.28 379.62 ;
   RECT 23.18 379.62 933.28 381.33 ;
   RECT 23.18 381.33 933.28 383.04 ;
   RECT 23.18 383.04 933.28 384.75 ;
   RECT 23.18 384.75 933.28 386.46 ;
   RECT 23.18 386.46 933.28 388.17 ;
   RECT 23.18 388.17 933.28 389.88 ;
   RECT 23.18 389.88 933.28 391.59 ;
   RECT 23.18 391.59 933.28 393.3 ;
   RECT 23.18 393.3 933.28 395.01 ;
   RECT 23.18 395.01 933.28 396.72 ;
   RECT 23.18 396.72 933.28 398.43 ;
   RECT 23.18 398.43 933.28 400.14 ;
   RECT 23.18 400.14 933.28 401.85 ;
   RECT 23.18 401.85 933.28 403.56 ;
   RECT 23.18 403.56 933.28 405.27 ;
   RECT 23.18 405.27 933.28 406.98 ;
   RECT 23.18 406.98 933.28 408.69 ;
   RECT 23.18 408.69 933.28 410.4 ;
   RECT 23.18 410.4 933.28 412.11 ;
   RECT 23.18 412.11 933.28 413.82 ;
   RECT 23.18 413.82 933.28 415.53 ;
   RECT 23.18 415.53 933.28 417.24 ;
   RECT 23.18 417.24 933.28 418.95 ;
   RECT 23.18 418.95 933.28 420.66 ;
   RECT 23.18 420.66 933.28 422.37 ;
   RECT 23.18 422.37 933.28 424.08 ;
   RECT 23.18 424.08 933.28 425.79 ;
   RECT 23.18 425.79 933.28 427.5 ;
   RECT 23.18 427.5 933.28 429.21 ;
   RECT 23.18 429.21 933.28 430.92 ;
   RECT 0.0 430.92 933.28 432.63 ;
   RECT 0.0 432.63 933.28 434.34 ;
   RECT 0.0 434.34 933.28 436.05 ;
   RECT 0.0 436.05 933.28 437.76 ;
   RECT 0.0 437.76 933.28 439.47 ;
   RECT 0.0 439.47 933.28 441.18 ;
   RECT 0.0 441.18 933.28 442.89 ;
   RECT 0.0 442.89 933.28 444.6 ;
   RECT 0.0 444.6 933.28 446.31 ;
   RECT 0.0 446.31 933.28 448.02 ;
   RECT 0.0 448.02 933.28 449.73 ;
   RECT 0.0 449.73 933.28 451.44 ;
   RECT 0.0 451.44 933.28 453.15 ;
   RECT 0.0 453.15 933.28 454.86 ;
   RECT 0.0 454.86 933.28 456.57 ;
   RECT 0.0 456.57 933.28 458.28 ;
   RECT 0.0 458.28 933.28 459.99 ;
   RECT 23.18 459.99 933.28 461.7 ;
   RECT 23.18 461.7 933.28 463.41 ;
   RECT 23.18 463.41 933.28 465.12 ;
   RECT 23.18 465.12 933.28 466.83 ;
   RECT 23.18 466.83 933.28 468.54 ;
   RECT 23.18 468.54 933.28 470.25 ;
   RECT 23.18 470.25 933.28 471.96 ;
   RECT 23.18 471.96 933.28 473.67 ;
   RECT 23.18 473.67 933.28 475.38 ;
   RECT 23.18 475.38 933.28 477.09 ;
   RECT 23.18 477.09 933.28 478.8 ;
   RECT 23.18 478.8 933.28 480.51 ;
   RECT 23.18 480.51 933.28 482.22 ;
   RECT 23.18 482.22 933.28 483.93 ;
   RECT 23.18 483.93 933.28 485.64 ;
   RECT 23.18 485.64 933.28 487.35 ;
   RECT 23.18 487.35 933.28 489.06 ;
   RECT 23.18 489.06 933.28 490.77 ;
   RECT 23.18 490.77 933.28 492.48 ;
   RECT 23.18 492.48 933.28 494.19 ;
   RECT 23.18 494.19 933.28 495.9 ;
   RECT 23.18 495.9 933.28 497.61 ;
   RECT 23.18 497.61 933.28 499.32 ;
   RECT 23.18 499.32 933.28 501.03 ;
   RECT 23.18 501.03 933.28 502.74 ;
   RECT 23.18 502.74 933.28 504.45 ;
   RECT 23.18 504.45 933.28 506.16 ;
   RECT 23.18 506.16 933.28 507.87 ;
   RECT 23.18 507.87 933.28 509.58 ;
   RECT 23.18 509.58 933.28 511.29 ;
   RECT 23.18 511.29 933.28 513.0 ;
   RECT 23.18 513.0 933.28 514.71 ;
   RECT 23.18 514.71 933.28 516.42 ;
   RECT 23.18 516.42 933.28 518.13 ;
   RECT 23.18 518.13 933.28 519.84 ;
   RECT 23.18 519.84 933.28 521.55 ;
   RECT 23.18 521.55 933.28 523.26 ;
   RECT 23.18 523.26 933.28 524.97 ;
   RECT 23.18 524.97 933.28 526.68 ;
   RECT 23.18 526.68 933.28 528.39 ;
   RECT 23.18 528.39 933.28 530.1 ;
   RECT 23.18 530.1 933.28 531.81 ;
   RECT 23.18 531.81 933.28 533.52 ;
   RECT 23.18 533.52 933.28 535.23 ;
   RECT 23.18 535.23 933.28 536.94 ;
   RECT 23.18 536.94 933.28 538.65 ;
   RECT 23.18 538.65 933.28 540.36 ;
   RECT 23.18 540.36 933.28 542.07 ;
   RECT 23.18 542.07 933.28 543.78 ;
   RECT 23.18 543.78 933.28 545.49 ;
   RECT 23.18 545.49 933.28 547.2 ;
   RECT 23.18 547.2 933.28 548.91 ;
   RECT 23.18 548.91 933.28 550.62 ;
   RECT 23.18 550.62 933.28 552.33 ;
   RECT 23.18 552.33 933.28 554.04 ;
   RECT 23.18 554.04 933.28 555.75 ;
   RECT 23.18 555.75 933.28 557.46 ;
   RECT 23.18 557.46 933.28 559.17 ;
   RECT 23.18 559.17 933.28 560.88 ;
   RECT 23.18 560.88 933.28 562.59 ;
   RECT 23.18 562.59 933.28 564.3 ;
   RECT 23.18 564.3 933.28 566.01 ;
   RECT 23.18 566.01 933.28 567.72 ;
   RECT 23.18 567.72 933.28 569.43 ;
   RECT 23.18 569.43 933.28 571.14 ;
   RECT 23.18 571.14 933.28 572.85 ;
   RECT 23.18 572.85 933.28 574.56 ;
   RECT 23.18 574.56 933.28 576.27 ;
   RECT 23.18 576.27 933.28 577.98 ;
   RECT 23.18 577.98 933.28 579.69 ;
   RECT 23.18 579.69 933.28 581.4 ;
   RECT 23.18 581.4 933.28 583.11 ;
   RECT 23.18 583.11 933.28 584.82 ;
   RECT 23.18 584.82 933.28 586.53 ;
   RECT 23.18 586.53 933.28 588.24 ;
   RECT 23.18 588.24 933.28 589.95 ;
   RECT 23.18 589.95 933.28 591.66 ;
   RECT 23.18 591.66 933.28 593.37 ;
   RECT 23.18 593.37 933.28 595.08 ;
   RECT 23.18 595.08 933.28 596.79 ;
   RECT 23.18 596.79 933.28 598.5 ;
   RECT 23.18 598.5 933.28 600.21 ;
   RECT 23.18 600.21 933.28 601.92 ;
   RECT 23.18 601.92 933.28 603.63 ;
   RECT 23.18 603.63 933.28 605.34 ;
   RECT 23.18 605.34 933.28 607.05 ;
   RECT 23.18 607.05 933.28 608.76 ;
   RECT 23.18 608.76 933.28 610.47 ;
   RECT 23.18 610.47 933.28 612.18 ;
   RECT 23.18 612.18 933.28 613.89 ;
   RECT 23.18 613.89 933.28 615.6 ;
   RECT 23.18 615.6 933.28 617.31 ;
   RECT 23.18 617.31 933.28 619.02 ;
   RECT 23.18 619.02 933.28 620.73 ;
   RECT 23.18 620.73 933.28 622.44 ;
   RECT 23.18 622.44 933.28 624.15 ;
   RECT 23.18 624.15 933.28 625.86 ;
   RECT 23.18 625.86 933.28 627.57 ;
   RECT 23.18 627.57 933.28 629.28 ;
   RECT 23.18 629.28 933.28 630.99 ;
   RECT 23.18 630.99 933.28 632.7 ;
   RECT 23.18 632.7 933.28 634.41 ;
   RECT 23.18 634.41 933.28 636.12 ;
   RECT 23.18 636.12 933.28 637.83 ;
   RECT 23.18 637.83 933.28 639.54 ;
   RECT 23.18 639.54 933.28 641.25 ;
   RECT 23.18 641.25 933.28 642.96 ;
   RECT 23.18 642.96 933.28 644.67 ;
   RECT 23.18 644.67 933.28 646.38 ;
   RECT 23.18 646.38 933.28 648.09 ;
   RECT 23.18 648.09 933.28 649.8 ;
   RECT 23.18 649.8 933.28 651.51 ;
   RECT 23.18 651.51 933.28 653.22 ;
   RECT 23.18 653.22 933.28 654.93 ;
   RECT 23.18 654.93 933.28 656.64 ;
   RECT 23.18 656.64 933.28 658.35 ;
   RECT 23.18 658.35 933.28 660.06 ;
   RECT 23.18 660.06 933.28 661.77 ;
   RECT 23.18 661.77 933.28 663.48 ;
   RECT 23.18 663.48 933.28 665.19 ;
   RECT 23.18 665.19 933.28 666.9 ;
   RECT 23.18 666.9 933.28 668.61 ;
   RECT 23.18 668.61 933.28 670.32 ;
   RECT 23.18 670.32 933.28 672.03 ;
   RECT 23.18 672.03 933.28 673.74 ;
   RECT 23.18 673.74 933.28 675.45 ;
   RECT 23.18 675.45 933.28 677.16 ;
   RECT 23.18 677.16 933.28 678.87 ;
   RECT 23.18 678.87 933.28 680.58 ;
   RECT 23.18 680.58 933.28 682.29 ;
   RECT 23.18 682.29 933.28 684.0 ;
   RECT 23.18 684.0 933.28 685.71 ;
   RECT 23.18 685.71 933.28 687.42 ;
   RECT 23.18 687.42 933.28 689.13 ;
   RECT 23.18 689.13 933.28 690.84 ;
   RECT 23.18 690.84 933.28 692.55 ;
   RECT 23.18 692.55 933.28 694.26 ;
   RECT 23.18 694.26 933.28 695.97 ;
   RECT 23.18 695.97 933.28 697.68 ;
   RECT 23.18 697.68 933.28 699.39 ;
   RECT 23.18 699.39 933.28 701.1 ;
   RECT 23.18 701.1 933.28 702.81 ;
   RECT 23.18 702.81 933.28 704.52 ;
   RECT 23.18 704.52 933.28 706.23 ;
   RECT 23.18 706.23 933.28 707.94 ;
   RECT 23.18 707.94 933.28 709.65 ;
   RECT 23.18 709.65 933.28 711.36 ;
   RECT 23.18 711.36 933.28 713.07 ;
   RECT 23.18 713.07 933.28 714.78 ;
   RECT 23.18 714.78 933.28 716.49 ;
   RECT 23.18 716.49 933.28 718.2 ;
   RECT 23.18 718.2 933.28 719.91 ;
   RECT 23.18 719.91 933.28 721.62 ;
   RECT 23.18 721.62 933.28 723.33 ;
   RECT 23.18 723.33 933.28 725.04 ;
   RECT 23.18 725.04 933.28 726.75 ;
   RECT 23.18 726.75 933.28 728.46 ;
   RECT 23.18 728.46 933.28 730.17 ;
   RECT 23.18 730.17 933.28 731.88 ;
   RECT 23.18 731.88 933.28 733.59 ;
   RECT 23.18 733.59 933.28 735.3 ;
   RECT 23.18 735.3 933.28 737.01 ;
   RECT 23.18 737.01 933.28 738.72 ;
   RECT 23.18 738.72 933.28 740.43 ;
   RECT 23.18 740.43 933.28 742.14 ;
   RECT 23.18 742.14 933.28 743.85 ;
   RECT 23.18 743.85 933.28 745.56 ;
   RECT 23.18 745.56 933.28 747.27 ;
   RECT 23.18 747.27 933.28 748.98 ;
   RECT 23.18 748.98 933.28 750.69 ;
   RECT 23.18 750.69 933.28 752.4 ;
   RECT 23.18 752.4 933.28 754.11 ;
   RECT 23.18 754.11 933.28 755.82 ;
   RECT 23.18 755.82 933.28 757.53 ;
   RECT 23.18 757.53 933.28 759.24 ;
   RECT 23.18 759.24 933.28 760.95 ;
   RECT 23.18 760.95 933.28 762.66 ;
   RECT 23.18 762.66 933.28 764.37 ;
   RECT 23.18 764.37 933.28 766.08 ;
   RECT 23.18 766.08 933.28 767.79 ;
   RECT 23.18 767.79 933.28 769.5 ;
   RECT 23.18 769.5 933.28 771.21 ;
   RECT 23.18 771.21 933.28 772.92 ;
   RECT 23.18 772.92 933.28 774.63 ;
   RECT 23.18 774.63 933.28 776.34 ;
   RECT 23.18 776.34 933.28 778.05 ;
   RECT 23.18 778.05 933.28 779.76 ;
   RECT 23.18 779.76 933.28 781.47 ;
   RECT 23.18 781.47 933.28 783.18 ;
   RECT 23.18 783.18 933.28 784.89 ;
   RECT 23.18 784.89 933.28 786.6 ;
   RECT 23.18 786.6 933.28 788.31 ;
   RECT 23.18 788.31 933.28 790.02 ;
   RECT 23.18 790.02 933.28 791.73 ;
   RECT 23.18 791.73 933.28 793.44 ;
   RECT 23.18 793.44 933.28 795.15 ;
   RECT 23.18 795.15 933.28 796.86 ;
   RECT 23.18 796.86 933.28 798.57 ;
   RECT 23.18 798.57 933.28 800.28 ;
   RECT 23.18 800.28 933.28 801.99 ;
   RECT 23.18 801.99 933.28 803.7 ;
   RECT 23.18 803.7 933.28 805.41 ;
   RECT 23.18 805.41 933.28 807.12 ;
   RECT 23.18 807.12 933.28 808.83 ;
   RECT 23.18 808.83 933.28 810.54 ;
   RECT 23.18 810.54 933.28 812.25 ;
   RECT 23.18 812.25 933.28 813.96 ;
   RECT 23.18 813.96 933.28 815.67 ;
   RECT 23.18 815.67 933.28 817.38 ;
   RECT 23.18 817.38 933.28 819.09 ;
   RECT 23.18 819.09 933.28 820.8 ;
   RECT 23.18 820.8 933.28 822.51 ;
   RECT 23.18 822.51 933.28 824.22 ;
   RECT 23.18 824.22 933.28 825.93 ;
   RECT 23.18 825.93 933.28 827.64 ;
   RECT 23.18 827.64 933.28 829.35 ;
   RECT 23.18 829.35 933.28 831.06 ;
   RECT 23.18 831.06 933.28 832.77 ;
   RECT 23.18 832.77 933.28 834.48 ;
   RECT 23.18 834.48 933.28 836.19 ;
   RECT 23.18 836.19 933.28 837.9 ;
   RECT 23.18 837.9 933.28 839.61 ;
   RECT 23.18 839.61 933.28 841.32 ;
   RECT 23.18 841.32 933.28 843.03 ;
   RECT 23.18 843.03 933.28 844.74 ;
   RECT 23.18 844.74 933.28 846.45 ;
   RECT 23.18 846.45 933.28 848.16 ;
   RECT 23.18 848.16 933.28 849.87 ;
   RECT 23.18 849.87 933.28 851.58 ;
   RECT 23.18 851.58 933.28 853.29 ;
   RECT 23.18 853.29 933.28 855.0 ;
   RECT 23.18 855.0 933.28 856.71 ;
   RECT 23.18 856.71 933.28 858.42 ;
   RECT 23.18 858.42 933.28 860.13 ;
   RECT 23.18 860.13 933.28 861.84 ;
   RECT 23.18 861.84 933.28 863.55 ;
   RECT 23.18 863.55 933.28 865.26 ;
   RECT 23.18 865.26 933.28 866.97 ;
   RECT 23.18 866.97 933.28 868.68 ;
   RECT 23.18 868.68 933.28 870.39 ;
   RECT 23.18 870.39 933.28 872.1 ;
   RECT 23.18 872.1 933.28 873.81 ;
   RECT 23.18 873.81 933.28 875.52 ;
   RECT 23.18 875.52 933.28 877.23 ;
   RECT 23.18 877.23 933.28 878.94 ;
  LAYER via1 ;
   RECT 23.18 0.0 933.28 1.71 ;
   RECT 23.18 1.71 933.28 3.42 ;
   RECT 23.18 3.42 933.28 5.13 ;
   RECT 23.18 5.13 933.28 6.84 ;
   RECT 23.18 6.84 933.28 8.55 ;
   RECT 23.18 8.55 933.28 10.26 ;
   RECT 23.18 10.26 933.28 11.97 ;
   RECT 23.18 11.97 933.28 13.68 ;
   RECT 23.18 13.68 933.28 15.39 ;
   RECT 23.18 15.39 933.28 17.1 ;
   RECT 23.18 17.1 933.28 18.81 ;
   RECT 23.18 18.81 933.28 20.52 ;
   RECT 23.18 20.52 933.28 22.23 ;
   RECT 23.18 22.23 933.28 23.94 ;
   RECT 23.18 23.94 933.28 25.65 ;
   RECT 23.18 25.65 933.28 27.36 ;
   RECT 23.18 27.36 933.28 29.07 ;
   RECT 23.18 29.07 933.28 30.78 ;
   RECT 23.18 30.78 933.28 32.49 ;
   RECT 23.18 32.49 933.28 34.2 ;
   RECT 23.18 34.2 933.28 35.91 ;
   RECT 23.18 35.91 933.28 37.62 ;
   RECT 23.18 37.62 933.28 39.33 ;
   RECT 23.18 39.33 933.28 41.04 ;
   RECT 23.18 41.04 933.28 42.75 ;
   RECT 23.18 42.75 933.28 44.46 ;
   RECT 23.18 44.46 933.28 46.17 ;
   RECT 23.18 46.17 933.28 47.88 ;
   RECT 23.18 47.88 933.28 49.59 ;
   RECT 23.18 49.59 933.28 51.3 ;
   RECT 23.18 51.3 933.28 53.01 ;
   RECT 23.18 53.01 933.28 54.72 ;
   RECT 23.18 54.72 933.28 56.43 ;
   RECT 23.18 56.43 933.28 58.14 ;
   RECT 23.18 58.14 933.28 59.85 ;
   RECT 23.18 59.85 933.28 61.56 ;
   RECT 23.18 61.56 933.28 63.27 ;
   RECT 23.18 63.27 933.28 64.98 ;
   RECT 23.18 64.98 933.28 66.69 ;
   RECT 23.18 66.69 933.28 68.4 ;
   RECT 23.18 68.4 933.28 70.11 ;
   RECT 23.18 70.11 933.28 71.82 ;
   RECT 23.18 71.82 933.28 73.53 ;
   RECT 23.18 73.53 933.28 75.24 ;
   RECT 23.18 75.24 933.28 76.95 ;
   RECT 23.18 76.95 933.28 78.66 ;
   RECT 23.18 78.66 933.28 80.37 ;
   RECT 23.18 80.37 933.28 82.08 ;
   RECT 23.18 82.08 933.28 83.79 ;
   RECT 23.18 83.79 933.28 85.5 ;
   RECT 23.18 85.5 933.28 87.21 ;
   RECT 23.18 87.21 933.28 88.92 ;
   RECT 23.18 88.92 933.28 90.63 ;
   RECT 23.18 90.63 933.28 92.34 ;
   RECT 23.18 92.34 933.28 94.05 ;
   RECT 23.18 94.05 933.28 95.76 ;
   RECT 23.18 95.76 933.28 97.47 ;
   RECT 23.18 97.47 933.28 99.18 ;
   RECT 23.18 99.18 933.28 100.89 ;
   RECT 23.18 100.89 933.28 102.6 ;
   RECT 23.18 102.6 933.28 104.31 ;
   RECT 23.18 104.31 933.28 106.02 ;
   RECT 23.18 106.02 933.28 107.73 ;
   RECT 23.18 107.73 933.28 109.44 ;
   RECT 23.18 109.44 933.28 111.15 ;
   RECT 23.18 111.15 933.28 112.86 ;
   RECT 23.18 112.86 933.28 114.57 ;
   RECT 23.18 114.57 933.28 116.28 ;
   RECT 23.18 116.28 933.28 117.99 ;
   RECT 23.18 117.99 933.28 119.7 ;
   RECT 23.18 119.7 933.28 121.41 ;
   RECT 23.18 121.41 933.28 123.12 ;
   RECT 23.18 123.12 933.28 124.83 ;
   RECT 23.18 124.83 933.28 126.54 ;
   RECT 23.18 126.54 933.28 128.25 ;
   RECT 23.18 128.25 933.28 129.96 ;
   RECT 23.18 129.96 933.28 131.67 ;
   RECT 23.18 131.67 933.28 133.38 ;
   RECT 23.18 133.38 933.28 135.09 ;
   RECT 23.18 135.09 933.28 136.8 ;
   RECT 23.18 136.8 933.28 138.51 ;
   RECT 23.18 138.51 933.28 140.22 ;
   RECT 23.18 140.22 933.28 141.93 ;
   RECT 23.18 141.93 933.28 143.64 ;
   RECT 23.18 143.64 933.28 145.35 ;
   RECT 23.18 145.35 933.28 147.06 ;
   RECT 23.18 147.06 933.28 148.77 ;
   RECT 23.18 148.77 933.28 150.48 ;
   RECT 23.18 150.48 933.28 152.19 ;
   RECT 23.18 152.19 933.28 153.9 ;
   RECT 23.18 153.9 933.28 155.61 ;
   RECT 23.18 155.61 933.28 157.32 ;
   RECT 23.18 157.32 933.28 159.03 ;
   RECT 23.18 159.03 933.28 160.74 ;
   RECT 23.18 160.74 933.28 162.45 ;
   RECT 23.18 162.45 933.28 164.16 ;
   RECT 23.18 164.16 933.28 165.87 ;
   RECT 23.18 165.87 933.28 167.58 ;
   RECT 23.18 167.58 933.28 169.29 ;
   RECT 23.18 169.29 933.28 171.0 ;
   RECT 23.18 171.0 933.28 172.71 ;
   RECT 23.18 172.71 933.28 174.42 ;
   RECT 23.18 174.42 933.28 176.13 ;
   RECT 23.18 176.13 933.28 177.84 ;
   RECT 23.18 177.84 933.28 179.55 ;
   RECT 23.18 179.55 933.28 181.26 ;
   RECT 23.18 181.26 933.28 182.97 ;
   RECT 23.18 182.97 933.28 184.68 ;
   RECT 23.18 184.68 933.28 186.39 ;
   RECT 23.18 186.39 933.28 188.1 ;
   RECT 23.18 188.1 933.28 189.81 ;
   RECT 23.18 189.81 933.28 191.52 ;
   RECT 23.18 191.52 933.28 193.23 ;
   RECT 23.18 193.23 933.28 194.94 ;
   RECT 23.18 194.94 933.28 196.65 ;
   RECT 23.18 196.65 933.28 198.36 ;
   RECT 23.18 198.36 933.28 200.07 ;
   RECT 23.18 200.07 933.28 201.78 ;
   RECT 23.18 201.78 933.28 203.49 ;
   RECT 23.18 203.49 933.28 205.2 ;
   RECT 23.18 205.2 933.28 206.91 ;
   RECT 23.18 206.91 933.28 208.62 ;
   RECT 23.18 208.62 933.28 210.33 ;
   RECT 23.18 210.33 933.28 212.04 ;
   RECT 23.18 212.04 933.28 213.75 ;
   RECT 23.18 213.75 933.28 215.46 ;
   RECT 23.18 215.46 933.28 217.17 ;
   RECT 23.18 217.17 933.28 218.88 ;
   RECT 23.18 218.88 933.28 220.59 ;
   RECT 23.18 220.59 933.28 222.3 ;
   RECT 23.18 222.3 933.28 224.01 ;
   RECT 23.18 224.01 933.28 225.72 ;
   RECT 23.18 225.72 933.28 227.43 ;
   RECT 23.18 227.43 933.28 229.14 ;
   RECT 23.18 229.14 933.28 230.85 ;
   RECT 23.18 230.85 933.28 232.56 ;
   RECT 23.18 232.56 933.28 234.27 ;
   RECT 23.18 234.27 933.28 235.98 ;
   RECT 23.18 235.98 933.28 237.69 ;
   RECT 23.18 237.69 933.28 239.4 ;
   RECT 23.18 239.4 933.28 241.11 ;
   RECT 23.18 241.11 933.28 242.82 ;
   RECT 23.18 242.82 933.28 244.53 ;
   RECT 23.18 244.53 933.28 246.24 ;
   RECT 23.18 246.24 933.28 247.95 ;
   RECT 23.18 247.95 933.28 249.66 ;
   RECT 23.18 249.66 933.28 251.37 ;
   RECT 23.18 251.37 933.28 253.08 ;
   RECT 23.18 253.08 933.28 254.79 ;
   RECT 23.18 254.79 933.28 256.5 ;
   RECT 23.18 256.5 933.28 258.21 ;
   RECT 23.18 258.21 933.28 259.92 ;
   RECT 23.18 259.92 933.28 261.63 ;
   RECT 23.18 261.63 933.28 263.34 ;
   RECT 23.18 263.34 933.28 265.05 ;
   RECT 23.18 265.05 933.28 266.76 ;
   RECT 23.18 266.76 933.28 268.47 ;
   RECT 23.18 268.47 933.28 270.18 ;
   RECT 23.18 270.18 933.28 271.89 ;
   RECT 23.18 271.89 933.28 273.6 ;
   RECT 23.18 273.6 933.28 275.31 ;
   RECT 23.18 275.31 933.28 277.02 ;
   RECT 23.18 277.02 933.28 278.73 ;
   RECT 23.18 278.73 933.28 280.44 ;
   RECT 23.18 280.44 933.28 282.15 ;
   RECT 23.18 282.15 933.28 283.86 ;
   RECT 23.18 283.86 933.28 285.57 ;
   RECT 23.18 285.57 933.28 287.28 ;
   RECT 23.18 287.28 933.28 288.99 ;
   RECT 23.18 288.99 933.28 290.7 ;
   RECT 23.18 290.7 933.28 292.41 ;
   RECT 23.18 292.41 933.28 294.12 ;
   RECT 23.18 294.12 933.28 295.83 ;
   RECT 23.18 295.83 933.28 297.54 ;
   RECT 23.18 297.54 933.28 299.25 ;
   RECT 23.18 299.25 933.28 300.96 ;
   RECT 23.18 300.96 933.28 302.67 ;
   RECT 23.18 302.67 933.28 304.38 ;
   RECT 23.18 304.38 933.28 306.09 ;
   RECT 23.18 306.09 933.28 307.8 ;
   RECT 23.18 307.8 933.28 309.51 ;
   RECT 23.18 309.51 933.28 311.22 ;
   RECT 23.18 311.22 933.28 312.93 ;
   RECT 23.18 312.93 933.28 314.64 ;
   RECT 23.18 314.64 933.28 316.35 ;
   RECT 23.18 316.35 933.28 318.06 ;
   RECT 23.18 318.06 933.28 319.77 ;
   RECT 23.18 319.77 933.28 321.48 ;
   RECT 23.18 321.48 933.28 323.19 ;
   RECT 23.18 323.19 933.28 324.9 ;
   RECT 23.18 324.9 933.28 326.61 ;
   RECT 23.18 326.61 933.28 328.32 ;
   RECT 23.18 328.32 933.28 330.03 ;
   RECT 23.18 330.03 933.28 331.74 ;
   RECT 23.18 331.74 933.28 333.45 ;
   RECT 23.18 333.45 933.28 335.16 ;
   RECT 23.18 335.16 933.28 336.87 ;
   RECT 23.18 336.87 933.28 338.58 ;
   RECT 23.18 338.58 933.28 340.29 ;
   RECT 23.18 340.29 933.28 342.0 ;
   RECT 23.18 342.0 933.28 343.71 ;
   RECT 23.18 343.71 933.28 345.42 ;
   RECT 23.18 345.42 933.28 347.13 ;
   RECT 23.18 347.13 933.28 348.84 ;
   RECT 23.18 348.84 933.28 350.55 ;
   RECT 23.18 350.55 933.28 352.26 ;
   RECT 23.18 352.26 933.28 353.97 ;
   RECT 23.18 353.97 933.28 355.68 ;
   RECT 23.18 355.68 933.28 357.39 ;
   RECT 23.18 357.39 933.28 359.1 ;
   RECT 23.18 359.1 933.28 360.81 ;
   RECT 23.18 360.81 933.28 362.52 ;
   RECT 23.18 362.52 933.28 364.23 ;
   RECT 23.18 364.23 933.28 365.94 ;
   RECT 23.18 365.94 933.28 367.65 ;
   RECT 23.18 367.65 933.28 369.36 ;
   RECT 23.18 369.36 933.28 371.07 ;
   RECT 23.18 371.07 933.28 372.78 ;
   RECT 23.18 372.78 933.28 374.49 ;
   RECT 23.18 374.49 933.28 376.2 ;
   RECT 23.18 376.2 933.28 377.91 ;
   RECT 23.18 377.91 933.28 379.62 ;
   RECT 23.18 379.62 933.28 381.33 ;
   RECT 23.18 381.33 933.28 383.04 ;
   RECT 23.18 383.04 933.28 384.75 ;
   RECT 23.18 384.75 933.28 386.46 ;
   RECT 23.18 386.46 933.28 388.17 ;
   RECT 23.18 388.17 933.28 389.88 ;
   RECT 23.18 389.88 933.28 391.59 ;
   RECT 23.18 391.59 933.28 393.3 ;
   RECT 23.18 393.3 933.28 395.01 ;
   RECT 23.18 395.01 933.28 396.72 ;
   RECT 23.18 396.72 933.28 398.43 ;
   RECT 23.18 398.43 933.28 400.14 ;
   RECT 23.18 400.14 933.28 401.85 ;
   RECT 23.18 401.85 933.28 403.56 ;
   RECT 23.18 403.56 933.28 405.27 ;
   RECT 23.18 405.27 933.28 406.98 ;
   RECT 23.18 406.98 933.28 408.69 ;
   RECT 23.18 408.69 933.28 410.4 ;
   RECT 23.18 410.4 933.28 412.11 ;
   RECT 23.18 412.11 933.28 413.82 ;
   RECT 23.18 413.82 933.28 415.53 ;
   RECT 23.18 415.53 933.28 417.24 ;
   RECT 23.18 417.24 933.28 418.95 ;
   RECT 23.18 418.95 933.28 420.66 ;
   RECT 23.18 420.66 933.28 422.37 ;
   RECT 23.18 422.37 933.28 424.08 ;
   RECT 23.18 424.08 933.28 425.79 ;
   RECT 23.18 425.79 933.28 427.5 ;
   RECT 23.18 427.5 933.28 429.21 ;
   RECT 23.18 429.21 933.28 430.92 ;
   RECT 0.0 430.92 933.28 432.63 ;
   RECT 0.0 432.63 933.28 434.34 ;
   RECT 0.0 434.34 933.28 436.05 ;
   RECT 0.0 436.05 933.28 437.76 ;
   RECT 0.0 437.76 933.28 439.47 ;
   RECT 0.0 439.47 933.28 441.18 ;
   RECT 0.0 441.18 933.28 442.89 ;
   RECT 0.0 442.89 933.28 444.6 ;
   RECT 0.0 444.6 933.28 446.31 ;
   RECT 0.0 446.31 933.28 448.02 ;
   RECT 0.0 448.02 933.28 449.73 ;
   RECT 0.0 449.73 933.28 451.44 ;
   RECT 0.0 451.44 933.28 453.15 ;
   RECT 0.0 453.15 933.28 454.86 ;
   RECT 0.0 454.86 933.28 456.57 ;
   RECT 0.0 456.57 933.28 458.28 ;
   RECT 0.0 458.28 933.28 459.99 ;
   RECT 23.18 459.99 933.28 461.7 ;
   RECT 23.18 461.7 933.28 463.41 ;
   RECT 23.18 463.41 933.28 465.12 ;
   RECT 23.18 465.12 933.28 466.83 ;
   RECT 23.18 466.83 933.28 468.54 ;
   RECT 23.18 468.54 933.28 470.25 ;
   RECT 23.18 470.25 933.28 471.96 ;
   RECT 23.18 471.96 933.28 473.67 ;
   RECT 23.18 473.67 933.28 475.38 ;
   RECT 23.18 475.38 933.28 477.09 ;
   RECT 23.18 477.09 933.28 478.8 ;
   RECT 23.18 478.8 933.28 480.51 ;
   RECT 23.18 480.51 933.28 482.22 ;
   RECT 23.18 482.22 933.28 483.93 ;
   RECT 23.18 483.93 933.28 485.64 ;
   RECT 23.18 485.64 933.28 487.35 ;
   RECT 23.18 487.35 933.28 489.06 ;
   RECT 23.18 489.06 933.28 490.77 ;
   RECT 23.18 490.77 933.28 492.48 ;
   RECT 23.18 492.48 933.28 494.19 ;
   RECT 23.18 494.19 933.28 495.9 ;
   RECT 23.18 495.9 933.28 497.61 ;
   RECT 23.18 497.61 933.28 499.32 ;
   RECT 23.18 499.32 933.28 501.03 ;
   RECT 23.18 501.03 933.28 502.74 ;
   RECT 23.18 502.74 933.28 504.45 ;
   RECT 23.18 504.45 933.28 506.16 ;
   RECT 23.18 506.16 933.28 507.87 ;
   RECT 23.18 507.87 933.28 509.58 ;
   RECT 23.18 509.58 933.28 511.29 ;
   RECT 23.18 511.29 933.28 513.0 ;
   RECT 23.18 513.0 933.28 514.71 ;
   RECT 23.18 514.71 933.28 516.42 ;
   RECT 23.18 516.42 933.28 518.13 ;
   RECT 23.18 518.13 933.28 519.84 ;
   RECT 23.18 519.84 933.28 521.55 ;
   RECT 23.18 521.55 933.28 523.26 ;
   RECT 23.18 523.26 933.28 524.97 ;
   RECT 23.18 524.97 933.28 526.68 ;
   RECT 23.18 526.68 933.28 528.39 ;
   RECT 23.18 528.39 933.28 530.1 ;
   RECT 23.18 530.1 933.28 531.81 ;
   RECT 23.18 531.81 933.28 533.52 ;
   RECT 23.18 533.52 933.28 535.23 ;
   RECT 23.18 535.23 933.28 536.94 ;
   RECT 23.18 536.94 933.28 538.65 ;
   RECT 23.18 538.65 933.28 540.36 ;
   RECT 23.18 540.36 933.28 542.07 ;
   RECT 23.18 542.07 933.28 543.78 ;
   RECT 23.18 543.78 933.28 545.49 ;
   RECT 23.18 545.49 933.28 547.2 ;
   RECT 23.18 547.2 933.28 548.91 ;
   RECT 23.18 548.91 933.28 550.62 ;
   RECT 23.18 550.62 933.28 552.33 ;
   RECT 23.18 552.33 933.28 554.04 ;
   RECT 23.18 554.04 933.28 555.75 ;
   RECT 23.18 555.75 933.28 557.46 ;
   RECT 23.18 557.46 933.28 559.17 ;
   RECT 23.18 559.17 933.28 560.88 ;
   RECT 23.18 560.88 933.28 562.59 ;
   RECT 23.18 562.59 933.28 564.3 ;
   RECT 23.18 564.3 933.28 566.01 ;
   RECT 23.18 566.01 933.28 567.72 ;
   RECT 23.18 567.72 933.28 569.43 ;
   RECT 23.18 569.43 933.28 571.14 ;
   RECT 23.18 571.14 933.28 572.85 ;
   RECT 23.18 572.85 933.28 574.56 ;
   RECT 23.18 574.56 933.28 576.27 ;
   RECT 23.18 576.27 933.28 577.98 ;
   RECT 23.18 577.98 933.28 579.69 ;
   RECT 23.18 579.69 933.28 581.4 ;
   RECT 23.18 581.4 933.28 583.11 ;
   RECT 23.18 583.11 933.28 584.82 ;
   RECT 23.18 584.82 933.28 586.53 ;
   RECT 23.18 586.53 933.28 588.24 ;
   RECT 23.18 588.24 933.28 589.95 ;
   RECT 23.18 589.95 933.28 591.66 ;
   RECT 23.18 591.66 933.28 593.37 ;
   RECT 23.18 593.37 933.28 595.08 ;
   RECT 23.18 595.08 933.28 596.79 ;
   RECT 23.18 596.79 933.28 598.5 ;
   RECT 23.18 598.5 933.28 600.21 ;
   RECT 23.18 600.21 933.28 601.92 ;
   RECT 23.18 601.92 933.28 603.63 ;
   RECT 23.18 603.63 933.28 605.34 ;
   RECT 23.18 605.34 933.28 607.05 ;
   RECT 23.18 607.05 933.28 608.76 ;
   RECT 23.18 608.76 933.28 610.47 ;
   RECT 23.18 610.47 933.28 612.18 ;
   RECT 23.18 612.18 933.28 613.89 ;
   RECT 23.18 613.89 933.28 615.6 ;
   RECT 23.18 615.6 933.28 617.31 ;
   RECT 23.18 617.31 933.28 619.02 ;
   RECT 23.18 619.02 933.28 620.73 ;
   RECT 23.18 620.73 933.28 622.44 ;
   RECT 23.18 622.44 933.28 624.15 ;
   RECT 23.18 624.15 933.28 625.86 ;
   RECT 23.18 625.86 933.28 627.57 ;
   RECT 23.18 627.57 933.28 629.28 ;
   RECT 23.18 629.28 933.28 630.99 ;
   RECT 23.18 630.99 933.28 632.7 ;
   RECT 23.18 632.7 933.28 634.41 ;
   RECT 23.18 634.41 933.28 636.12 ;
   RECT 23.18 636.12 933.28 637.83 ;
   RECT 23.18 637.83 933.28 639.54 ;
   RECT 23.18 639.54 933.28 641.25 ;
   RECT 23.18 641.25 933.28 642.96 ;
   RECT 23.18 642.96 933.28 644.67 ;
   RECT 23.18 644.67 933.28 646.38 ;
   RECT 23.18 646.38 933.28 648.09 ;
   RECT 23.18 648.09 933.28 649.8 ;
   RECT 23.18 649.8 933.28 651.51 ;
   RECT 23.18 651.51 933.28 653.22 ;
   RECT 23.18 653.22 933.28 654.93 ;
   RECT 23.18 654.93 933.28 656.64 ;
   RECT 23.18 656.64 933.28 658.35 ;
   RECT 23.18 658.35 933.28 660.06 ;
   RECT 23.18 660.06 933.28 661.77 ;
   RECT 23.18 661.77 933.28 663.48 ;
   RECT 23.18 663.48 933.28 665.19 ;
   RECT 23.18 665.19 933.28 666.9 ;
   RECT 23.18 666.9 933.28 668.61 ;
   RECT 23.18 668.61 933.28 670.32 ;
   RECT 23.18 670.32 933.28 672.03 ;
   RECT 23.18 672.03 933.28 673.74 ;
   RECT 23.18 673.74 933.28 675.45 ;
   RECT 23.18 675.45 933.28 677.16 ;
   RECT 23.18 677.16 933.28 678.87 ;
   RECT 23.18 678.87 933.28 680.58 ;
   RECT 23.18 680.58 933.28 682.29 ;
   RECT 23.18 682.29 933.28 684.0 ;
   RECT 23.18 684.0 933.28 685.71 ;
   RECT 23.18 685.71 933.28 687.42 ;
   RECT 23.18 687.42 933.28 689.13 ;
   RECT 23.18 689.13 933.28 690.84 ;
   RECT 23.18 690.84 933.28 692.55 ;
   RECT 23.18 692.55 933.28 694.26 ;
   RECT 23.18 694.26 933.28 695.97 ;
   RECT 23.18 695.97 933.28 697.68 ;
   RECT 23.18 697.68 933.28 699.39 ;
   RECT 23.18 699.39 933.28 701.1 ;
   RECT 23.18 701.1 933.28 702.81 ;
   RECT 23.18 702.81 933.28 704.52 ;
   RECT 23.18 704.52 933.28 706.23 ;
   RECT 23.18 706.23 933.28 707.94 ;
   RECT 23.18 707.94 933.28 709.65 ;
   RECT 23.18 709.65 933.28 711.36 ;
   RECT 23.18 711.36 933.28 713.07 ;
   RECT 23.18 713.07 933.28 714.78 ;
   RECT 23.18 714.78 933.28 716.49 ;
   RECT 23.18 716.49 933.28 718.2 ;
   RECT 23.18 718.2 933.28 719.91 ;
   RECT 23.18 719.91 933.28 721.62 ;
   RECT 23.18 721.62 933.28 723.33 ;
   RECT 23.18 723.33 933.28 725.04 ;
   RECT 23.18 725.04 933.28 726.75 ;
   RECT 23.18 726.75 933.28 728.46 ;
   RECT 23.18 728.46 933.28 730.17 ;
   RECT 23.18 730.17 933.28 731.88 ;
   RECT 23.18 731.88 933.28 733.59 ;
   RECT 23.18 733.59 933.28 735.3 ;
   RECT 23.18 735.3 933.28 737.01 ;
   RECT 23.18 737.01 933.28 738.72 ;
   RECT 23.18 738.72 933.28 740.43 ;
   RECT 23.18 740.43 933.28 742.14 ;
   RECT 23.18 742.14 933.28 743.85 ;
   RECT 23.18 743.85 933.28 745.56 ;
   RECT 23.18 745.56 933.28 747.27 ;
   RECT 23.18 747.27 933.28 748.98 ;
   RECT 23.18 748.98 933.28 750.69 ;
   RECT 23.18 750.69 933.28 752.4 ;
   RECT 23.18 752.4 933.28 754.11 ;
   RECT 23.18 754.11 933.28 755.82 ;
   RECT 23.18 755.82 933.28 757.53 ;
   RECT 23.18 757.53 933.28 759.24 ;
   RECT 23.18 759.24 933.28 760.95 ;
   RECT 23.18 760.95 933.28 762.66 ;
   RECT 23.18 762.66 933.28 764.37 ;
   RECT 23.18 764.37 933.28 766.08 ;
   RECT 23.18 766.08 933.28 767.79 ;
   RECT 23.18 767.79 933.28 769.5 ;
   RECT 23.18 769.5 933.28 771.21 ;
   RECT 23.18 771.21 933.28 772.92 ;
   RECT 23.18 772.92 933.28 774.63 ;
   RECT 23.18 774.63 933.28 776.34 ;
   RECT 23.18 776.34 933.28 778.05 ;
   RECT 23.18 778.05 933.28 779.76 ;
   RECT 23.18 779.76 933.28 781.47 ;
   RECT 23.18 781.47 933.28 783.18 ;
   RECT 23.18 783.18 933.28 784.89 ;
   RECT 23.18 784.89 933.28 786.6 ;
   RECT 23.18 786.6 933.28 788.31 ;
   RECT 23.18 788.31 933.28 790.02 ;
   RECT 23.18 790.02 933.28 791.73 ;
   RECT 23.18 791.73 933.28 793.44 ;
   RECT 23.18 793.44 933.28 795.15 ;
   RECT 23.18 795.15 933.28 796.86 ;
   RECT 23.18 796.86 933.28 798.57 ;
   RECT 23.18 798.57 933.28 800.28 ;
   RECT 23.18 800.28 933.28 801.99 ;
   RECT 23.18 801.99 933.28 803.7 ;
   RECT 23.18 803.7 933.28 805.41 ;
   RECT 23.18 805.41 933.28 807.12 ;
   RECT 23.18 807.12 933.28 808.83 ;
   RECT 23.18 808.83 933.28 810.54 ;
   RECT 23.18 810.54 933.28 812.25 ;
   RECT 23.18 812.25 933.28 813.96 ;
   RECT 23.18 813.96 933.28 815.67 ;
   RECT 23.18 815.67 933.28 817.38 ;
   RECT 23.18 817.38 933.28 819.09 ;
   RECT 23.18 819.09 933.28 820.8 ;
   RECT 23.18 820.8 933.28 822.51 ;
   RECT 23.18 822.51 933.28 824.22 ;
   RECT 23.18 824.22 933.28 825.93 ;
   RECT 23.18 825.93 933.28 827.64 ;
   RECT 23.18 827.64 933.28 829.35 ;
   RECT 23.18 829.35 933.28 831.06 ;
   RECT 23.18 831.06 933.28 832.77 ;
   RECT 23.18 832.77 933.28 834.48 ;
   RECT 23.18 834.48 933.28 836.19 ;
   RECT 23.18 836.19 933.28 837.9 ;
   RECT 23.18 837.9 933.28 839.61 ;
   RECT 23.18 839.61 933.28 841.32 ;
   RECT 23.18 841.32 933.28 843.03 ;
   RECT 23.18 843.03 933.28 844.74 ;
   RECT 23.18 844.74 933.28 846.45 ;
   RECT 23.18 846.45 933.28 848.16 ;
   RECT 23.18 848.16 933.28 849.87 ;
   RECT 23.18 849.87 933.28 851.58 ;
   RECT 23.18 851.58 933.28 853.29 ;
   RECT 23.18 853.29 933.28 855.0 ;
   RECT 23.18 855.0 933.28 856.71 ;
   RECT 23.18 856.71 933.28 858.42 ;
   RECT 23.18 858.42 933.28 860.13 ;
   RECT 23.18 860.13 933.28 861.84 ;
   RECT 23.18 861.84 933.28 863.55 ;
   RECT 23.18 863.55 933.28 865.26 ;
   RECT 23.18 865.26 933.28 866.97 ;
   RECT 23.18 866.97 933.28 868.68 ;
   RECT 23.18 868.68 933.28 870.39 ;
   RECT 23.18 870.39 933.28 872.1 ;
   RECT 23.18 872.1 933.28 873.81 ;
   RECT 23.18 873.81 933.28 875.52 ;
   RECT 23.18 875.52 933.28 877.23 ;
   RECT 23.18 877.23 933.28 878.94 ;
  LAYER metal2 ;
   RECT 23.18 0.0 933.28 1.71 ;
   RECT 23.18 1.71 933.28 3.42 ;
   RECT 23.18 3.42 933.28 5.13 ;
   RECT 23.18 5.13 933.28 6.84 ;
   RECT 23.18 6.84 933.28 8.55 ;
   RECT 23.18 8.55 933.28 10.26 ;
   RECT 23.18 10.26 933.28 11.97 ;
   RECT 23.18 11.97 933.28 13.68 ;
   RECT 23.18 13.68 933.28 15.39 ;
   RECT 23.18 15.39 933.28 17.1 ;
   RECT 23.18 17.1 933.28 18.81 ;
   RECT 23.18 18.81 933.28 20.52 ;
   RECT 23.18 20.52 933.28 22.23 ;
   RECT 23.18 22.23 933.28 23.94 ;
   RECT 23.18 23.94 933.28 25.65 ;
   RECT 23.18 25.65 933.28 27.36 ;
   RECT 23.18 27.36 933.28 29.07 ;
   RECT 23.18 29.07 933.28 30.78 ;
   RECT 23.18 30.78 933.28 32.49 ;
   RECT 23.18 32.49 933.28 34.2 ;
   RECT 23.18 34.2 933.28 35.91 ;
   RECT 23.18 35.91 933.28 37.62 ;
   RECT 23.18 37.62 933.28 39.33 ;
   RECT 23.18 39.33 933.28 41.04 ;
   RECT 23.18 41.04 933.28 42.75 ;
   RECT 23.18 42.75 933.28 44.46 ;
   RECT 23.18 44.46 933.28 46.17 ;
   RECT 23.18 46.17 933.28 47.88 ;
   RECT 23.18 47.88 933.28 49.59 ;
   RECT 23.18 49.59 933.28 51.3 ;
   RECT 23.18 51.3 933.28 53.01 ;
   RECT 23.18 53.01 933.28 54.72 ;
   RECT 23.18 54.72 933.28 56.43 ;
   RECT 23.18 56.43 933.28 58.14 ;
   RECT 23.18 58.14 933.28 59.85 ;
   RECT 23.18 59.85 933.28 61.56 ;
   RECT 23.18 61.56 933.28 63.27 ;
   RECT 23.18 63.27 933.28 64.98 ;
   RECT 23.18 64.98 933.28 66.69 ;
   RECT 23.18 66.69 933.28 68.4 ;
   RECT 23.18 68.4 933.28 70.11 ;
   RECT 23.18 70.11 933.28 71.82 ;
   RECT 23.18 71.82 933.28 73.53 ;
   RECT 23.18 73.53 933.28 75.24 ;
   RECT 23.18 75.24 933.28 76.95 ;
   RECT 23.18 76.95 933.28 78.66 ;
   RECT 23.18 78.66 933.28 80.37 ;
   RECT 23.18 80.37 933.28 82.08 ;
   RECT 23.18 82.08 933.28 83.79 ;
   RECT 23.18 83.79 933.28 85.5 ;
   RECT 23.18 85.5 933.28 87.21 ;
   RECT 23.18 87.21 933.28 88.92 ;
   RECT 23.18 88.92 933.28 90.63 ;
   RECT 23.18 90.63 933.28 92.34 ;
   RECT 23.18 92.34 933.28 94.05 ;
   RECT 23.18 94.05 933.28 95.76 ;
   RECT 23.18 95.76 933.28 97.47 ;
   RECT 23.18 97.47 933.28 99.18 ;
   RECT 23.18 99.18 933.28 100.89 ;
   RECT 23.18 100.89 933.28 102.6 ;
   RECT 23.18 102.6 933.28 104.31 ;
   RECT 23.18 104.31 933.28 106.02 ;
   RECT 23.18 106.02 933.28 107.73 ;
   RECT 23.18 107.73 933.28 109.44 ;
   RECT 23.18 109.44 933.28 111.15 ;
   RECT 23.18 111.15 933.28 112.86 ;
   RECT 23.18 112.86 933.28 114.57 ;
   RECT 23.18 114.57 933.28 116.28 ;
   RECT 23.18 116.28 933.28 117.99 ;
   RECT 23.18 117.99 933.28 119.7 ;
   RECT 23.18 119.7 933.28 121.41 ;
   RECT 23.18 121.41 933.28 123.12 ;
   RECT 23.18 123.12 933.28 124.83 ;
   RECT 23.18 124.83 933.28 126.54 ;
   RECT 23.18 126.54 933.28 128.25 ;
   RECT 23.18 128.25 933.28 129.96 ;
   RECT 23.18 129.96 933.28 131.67 ;
   RECT 23.18 131.67 933.28 133.38 ;
   RECT 23.18 133.38 933.28 135.09 ;
   RECT 23.18 135.09 933.28 136.8 ;
   RECT 23.18 136.8 933.28 138.51 ;
   RECT 23.18 138.51 933.28 140.22 ;
   RECT 23.18 140.22 933.28 141.93 ;
   RECT 23.18 141.93 933.28 143.64 ;
   RECT 23.18 143.64 933.28 145.35 ;
   RECT 23.18 145.35 933.28 147.06 ;
   RECT 23.18 147.06 933.28 148.77 ;
   RECT 23.18 148.77 933.28 150.48 ;
   RECT 23.18 150.48 933.28 152.19 ;
   RECT 23.18 152.19 933.28 153.9 ;
   RECT 23.18 153.9 933.28 155.61 ;
   RECT 23.18 155.61 933.28 157.32 ;
   RECT 23.18 157.32 933.28 159.03 ;
   RECT 23.18 159.03 933.28 160.74 ;
   RECT 23.18 160.74 933.28 162.45 ;
   RECT 23.18 162.45 933.28 164.16 ;
   RECT 23.18 164.16 933.28 165.87 ;
   RECT 23.18 165.87 933.28 167.58 ;
   RECT 23.18 167.58 933.28 169.29 ;
   RECT 23.18 169.29 933.28 171.0 ;
   RECT 23.18 171.0 933.28 172.71 ;
   RECT 23.18 172.71 933.28 174.42 ;
   RECT 23.18 174.42 933.28 176.13 ;
   RECT 23.18 176.13 933.28 177.84 ;
   RECT 23.18 177.84 933.28 179.55 ;
   RECT 23.18 179.55 933.28 181.26 ;
   RECT 23.18 181.26 933.28 182.97 ;
   RECT 23.18 182.97 933.28 184.68 ;
   RECT 23.18 184.68 933.28 186.39 ;
   RECT 23.18 186.39 933.28 188.1 ;
   RECT 23.18 188.1 933.28 189.81 ;
   RECT 23.18 189.81 933.28 191.52 ;
   RECT 23.18 191.52 933.28 193.23 ;
   RECT 23.18 193.23 933.28 194.94 ;
   RECT 23.18 194.94 933.28 196.65 ;
   RECT 23.18 196.65 933.28 198.36 ;
   RECT 23.18 198.36 933.28 200.07 ;
   RECT 23.18 200.07 933.28 201.78 ;
   RECT 23.18 201.78 933.28 203.49 ;
   RECT 23.18 203.49 933.28 205.2 ;
   RECT 23.18 205.2 933.28 206.91 ;
   RECT 23.18 206.91 933.28 208.62 ;
   RECT 23.18 208.62 933.28 210.33 ;
   RECT 23.18 210.33 933.28 212.04 ;
   RECT 23.18 212.04 933.28 213.75 ;
   RECT 23.18 213.75 933.28 215.46 ;
   RECT 23.18 215.46 933.28 217.17 ;
   RECT 23.18 217.17 933.28 218.88 ;
   RECT 23.18 218.88 933.28 220.59 ;
   RECT 23.18 220.59 933.28 222.3 ;
   RECT 23.18 222.3 933.28 224.01 ;
   RECT 23.18 224.01 933.28 225.72 ;
   RECT 23.18 225.72 933.28 227.43 ;
   RECT 23.18 227.43 933.28 229.14 ;
   RECT 23.18 229.14 933.28 230.85 ;
   RECT 23.18 230.85 933.28 232.56 ;
   RECT 23.18 232.56 933.28 234.27 ;
   RECT 23.18 234.27 933.28 235.98 ;
   RECT 23.18 235.98 933.28 237.69 ;
   RECT 23.18 237.69 933.28 239.4 ;
   RECT 23.18 239.4 933.28 241.11 ;
   RECT 23.18 241.11 933.28 242.82 ;
   RECT 23.18 242.82 933.28 244.53 ;
   RECT 23.18 244.53 933.28 246.24 ;
   RECT 23.18 246.24 933.28 247.95 ;
   RECT 23.18 247.95 933.28 249.66 ;
   RECT 23.18 249.66 933.28 251.37 ;
   RECT 23.18 251.37 933.28 253.08 ;
   RECT 23.18 253.08 933.28 254.79 ;
   RECT 23.18 254.79 933.28 256.5 ;
   RECT 23.18 256.5 933.28 258.21 ;
   RECT 23.18 258.21 933.28 259.92 ;
   RECT 23.18 259.92 933.28 261.63 ;
   RECT 23.18 261.63 933.28 263.34 ;
   RECT 23.18 263.34 933.28 265.05 ;
   RECT 23.18 265.05 933.28 266.76 ;
   RECT 23.18 266.76 933.28 268.47 ;
   RECT 23.18 268.47 933.28 270.18 ;
   RECT 23.18 270.18 933.28 271.89 ;
   RECT 23.18 271.89 933.28 273.6 ;
   RECT 23.18 273.6 933.28 275.31 ;
   RECT 23.18 275.31 933.28 277.02 ;
   RECT 23.18 277.02 933.28 278.73 ;
   RECT 23.18 278.73 933.28 280.44 ;
   RECT 23.18 280.44 933.28 282.15 ;
   RECT 23.18 282.15 933.28 283.86 ;
   RECT 23.18 283.86 933.28 285.57 ;
   RECT 23.18 285.57 933.28 287.28 ;
   RECT 23.18 287.28 933.28 288.99 ;
   RECT 23.18 288.99 933.28 290.7 ;
   RECT 23.18 290.7 933.28 292.41 ;
   RECT 23.18 292.41 933.28 294.12 ;
   RECT 23.18 294.12 933.28 295.83 ;
   RECT 23.18 295.83 933.28 297.54 ;
   RECT 23.18 297.54 933.28 299.25 ;
   RECT 23.18 299.25 933.28 300.96 ;
   RECT 23.18 300.96 933.28 302.67 ;
   RECT 23.18 302.67 933.28 304.38 ;
   RECT 23.18 304.38 933.28 306.09 ;
   RECT 23.18 306.09 933.28 307.8 ;
   RECT 23.18 307.8 933.28 309.51 ;
   RECT 23.18 309.51 933.28 311.22 ;
   RECT 23.18 311.22 933.28 312.93 ;
   RECT 23.18 312.93 933.28 314.64 ;
   RECT 23.18 314.64 933.28 316.35 ;
   RECT 23.18 316.35 933.28 318.06 ;
   RECT 23.18 318.06 933.28 319.77 ;
   RECT 23.18 319.77 933.28 321.48 ;
   RECT 23.18 321.48 933.28 323.19 ;
   RECT 23.18 323.19 933.28 324.9 ;
   RECT 23.18 324.9 933.28 326.61 ;
   RECT 23.18 326.61 933.28 328.32 ;
   RECT 23.18 328.32 933.28 330.03 ;
   RECT 23.18 330.03 933.28 331.74 ;
   RECT 23.18 331.74 933.28 333.45 ;
   RECT 23.18 333.45 933.28 335.16 ;
   RECT 23.18 335.16 933.28 336.87 ;
   RECT 23.18 336.87 933.28 338.58 ;
   RECT 23.18 338.58 933.28 340.29 ;
   RECT 23.18 340.29 933.28 342.0 ;
   RECT 23.18 342.0 933.28 343.71 ;
   RECT 23.18 343.71 933.28 345.42 ;
   RECT 23.18 345.42 933.28 347.13 ;
   RECT 23.18 347.13 933.28 348.84 ;
   RECT 23.18 348.84 933.28 350.55 ;
   RECT 23.18 350.55 933.28 352.26 ;
   RECT 23.18 352.26 933.28 353.97 ;
   RECT 23.18 353.97 933.28 355.68 ;
   RECT 23.18 355.68 933.28 357.39 ;
   RECT 23.18 357.39 933.28 359.1 ;
   RECT 23.18 359.1 933.28 360.81 ;
   RECT 23.18 360.81 933.28 362.52 ;
   RECT 23.18 362.52 933.28 364.23 ;
   RECT 23.18 364.23 933.28 365.94 ;
   RECT 23.18 365.94 933.28 367.65 ;
   RECT 23.18 367.65 933.28 369.36 ;
   RECT 23.18 369.36 933.28 371.07 ;
   RECT 23.18 371.07 933.28 372.78 ;
   RECT 23.18 372.78 933.28 374.49 ;
   RECT 23.18 374.49 933.28 376.2 ;
   RECT 23.18 376.2 933.28 377.91 ;
   RECT 23.18 377.91 933.28 379.62 ;
   RECT 23.18 379.62 933.28 381.33 ;
   RECT 23.18 381.33 933.28 383.04 ;
   RECT 23.18 383.04 933.28 384.75 ;
   RECT 23.18 384.75 933.28 386.46 ;
   RECT 23.18 386.46 933.28 388.17 ;
   RECT 23.18 388.17 933.28 389.88 ;
   RECT 23.18 389.88 933.28 391.59 ;
   RECT 23.18 391.59 933.28 393.3 ;
   RECT 23.18 393.3 933.28 395.01 ;
   RECT 23.18 395.01 933.28 396.72 ;
   RECT 23.18 396.72 933.28 398.43 ;
   RECT 23.18 398.43 933.28 400.14 ;
   RECT 23.18 400.14 933.28 401.85 ;
   RECT 23.18 401.85 933.28 403.56 ;
   RECT 23.18 403.56 933.28 405.27 ;
   RECT 23.18 405.27 933.28 406.98 ;
   RECT 23.18 406.98 933.28 408.69 ;
   RECT 23.18 408.69 933.28 410.4 ;
   RECT 23.18 410.4 933.28 412.11 ;
   RECT 23.18 412.11 933.28 413.82 ;
   RECT 23.18 413.82 933.28 415.53 ;
   RECT 23.18 415.53 933.28 417.24 ;
   RECT 23.18 417.24 933.28 418.95 ;
   RECT 23.18 418.95 933.28 420.66 ;
   RECT 23.18 420.66 933.28 422.37 ;
   RECT 23.18 422.37 933.28 424.08 ;
   RECT 23.18 424.08 933.28 425.79 ;
   RECT 23.18 425.79 933.28 427.5 ;
   RECT 23.18 427.5 933.28 429.21 ;
   RECT 23.18 429.21 933.28 430.92 ;
   RECT 0.0 430.92 933.28 432.63 ;
   RECT 0.0 432.63 933.28 434.34 ;
   RECT 0.0 434.34 933.28 436.05 ;
   RECT 0.0 436.05 933.28 437.76 ;
   RECT 0.0 437.76 933.28 439.47 ;
   RECT 0.0 439.47 933.28 441.18 ;
   RECT 0.0 441.18 933.28 442.89 ;
   RECT 0.0 442.89 933.28 444.6 ;
   RECT 0.0 444.6 933.28 446.31 ;
   RECT 0.0 446.31 933.28 448.02 ;
   RECT 0.0 448.02 933.28 449.73 ;
   RECT 0.0 449.73 933.28 451.44 ;
   RECT 0.0 451.44 933.28 453.15 ;
   RECT 0.0 453.15 933.28 454.86 ;
   RECT 0.0 454.86 933.28 456.57 ;
   RECT 0.0 456.57 933.28 458.28 ;
   RECT 0.0 458.28 933.28 459.99 ;
   RECT 23.18 459.99 933.28 461.7 ;
   RECT 23.18 461.7 933.28 463.41 ;
   RECT 23.18 463.41 933.28 465.12 ;
   RECT 23.18 465.12 933.28 466.83 ;
   RECT 23.18 466.83 933.28 468.54 ;
   RECT 23.18 468.54 933.28 470.25 ;
   RECT 23.18 470.25 933.28 471.96 ;
   RECT 23.18 471.96 933.28 473.67 ;
   RECT 23.18 473.67 933.28 475.38 ;
   RECT 23.18 475.38 933.28 477.09 ;
   RECT 23.18 477.09 933.28 478.8 ;
   RECT 23.18 478.8 933.28 480.51 ;
   RECT 23.18 480.51 933.28 482.22 ;
   RECT 23.18 482.22 933.28 483.93 ;
   RECT 23.18 483.93 933.28 485.64 ;
   RECT 23.18 485.64 933.28 487.35 ;
   RECT 23.18 487.35 933.28 489.06 ;
   RECT 23.18 489.06 933.28 490.77 ;
   RECT 23.18 490.77 933.28 492.48 ;
   RECT 23.18 492.48 933.28 494.19 ;
   RECT 23.18 494.19 933.28 495.9 ;
   RECT 23.18 495.9 933.28 497.61 ;
   RECT 23.18 497.61 933.28 499.32 ;
   RECT 23.18 499.32 933.28 501.03 ;
   RECT 23.18 501.03 933.28 502.74 ;
   RECT 23.18 502.74 933.28 504.45 ;
   RECT 23.18 504.45 933.28 506.16 ;
   RECT 23.18 506.16 933.28 507.87 ;
   RECT 23.18 507.87 933.28 509.58 ;
   RECT 23.18 509.58 933.28 511.29 ;
   RECT 23.18 511.29 933.28 513.0 ;
   RECT 23.18 513.0 933.28 514.71 ;
   RECT 23.18 514.71 933.28 516.42 ;
   RECT 23.18 516.42 933.28 518.13 ;
   RECT 23.18 518.13 933.28 519.84 ;
   RECT 23.18 519.84 933.28 521.55 ;
   RECT 23.18 521.55 933.28 523.26 ;
   RECT 23.18 523.26 933.28 524.97 ;
   RECT 23.18 524.97 933.28 526.68 ;
   RECT 23.18 526.68 933.28 528.39 ;
   RECT 23.18 528.39 933.28 530.1 ;
   RECT 23.18 530.1 933.28 531.81 ;
   RECT 23.18 531.81 933.28 533.52 ;
   RECT 23.18 533.52 933.28 535.23 ;
   RECT 23.18 535.23 933.28 536.94 ;
   RECT 23.18 536.94 933.28 538.65 ;
   RECT 23.18 538.65 933.28 540.36 ;
   RECT 23.18 540.36 933.28 542.07 ;
   RECT 23.18 542.07 933.28 543.78 ;
   RECT 23.18 543.78 933.28 545.49 ;
   RECT 23.18 545.49 933.28 547.2 ;
   RECT 23.18 547.2 933.28 548.91 ;
   RECT 23.18 548.91 933.28 550.62 ;
   RECT 23.18 550.62 933.28 552.33 ;
   RECT 23.18 552.33 933.28 554.04 ;
   RECT 23.18 554.04 933.28 555.75 ;
   RECT 23.18 555.75 933.28 557.46 ;
   RECT 23.18 557.46 933.28 559.17 ;
   RECT 23.18 559.17 933.28 560.88 ;
   RECT 23.18 560.88 933.28 562.59 ;
   RECT 23.18 562.59 933.28 564.3 ;
   RECT 23.18 564.3 933.28 566.01 ;
   RECT 23.18 566.01 933.28 567.72 ;
   RECT 23.18 567.72 933.28 569.43 ;
   RECT 23.18 569.43 933.28 571.14 ;
   RECT 23.18 571.14 933.28 572.85 ;
   RECT 23.18 572.85 933.28 574.56 ;
   RECT 23.18 574.56 933.28 576.27 ;
   RECT 23.18 576.27 933.28 577.98 ;
   RECT 23.18 577.98 933.28 579.69 ;
   RECT 23.18 579.69 933.28 581.4 ;
   RECT 23.18 581.4 933.28 583.11 ;
   RECT 23.18 583.11 933.28 584.82 ;
   RECT 23.18 584.82 933.28 586.53 ;
   RECT 23.18 586.53 933.28 588.24 ;
   RECT 23.18 588.24 933.28 589.95 ;
   RECT 23.18 589.95 933.28 591.66 ;
   RECT 23.18 591.66 933.28 593.37 ;
   RECT 23.18 593.37 933.28 595.08 ;
   RECT 23.18 595.08 933.28 596.79 ;
   RECT 23.18 596.79 933.28 598.5 ;
   RECT 23.18 598.5 933.28 600.21 ;
   RECT 23.18 600.21 933.28 601.92 ;
   RECT 23.18 601.92 933.28 603.63 ;
   RECT 23.18 603.63 933.28 605.34 ;
   RECT 23.18 605.34 933.28 607.05 ;
   RECT 23.18 607.05 933.28 608.76 ;
   RECT 23.18 608.76 933.28 610.47 ;
   RECT 23.18 610.47 933.28 612.18 ;
   RECT 23.18 612.18 933.28 613.89 ;
   RECT 23.18 613.89 933.28 615.6 ;
   RECT 23.18 615.6 933.28 617.31 ;
   RECT 23.18 617.31 933.28 619.02 ;
   RECT 23.18 619.02 933.28 620.73 ;
   RECT 23.18 620.73 933.28 622.44 ;
   RECT 23.18 622.44 933.28 624.15 ;
   RECT 23.18 624.15 933.28 625.86 ;
   RECT 23.18 625.86 933.28 627.57 ;
   RECT 23.18 627.57 933.28 629.28 ;
   RECT 23.18 629.28 933.28 630.99 ;
   RECT 23.18 630.99 933.28 632.7 ;
   RECT 23.18 632.7 933.28 634.41 ;
   RECT 23.18 634.41 933.28 636.12 ;
   RECT 23.18 636.12 933.28 637.83 ;
   RECT 23.18 637.83 933.28 639.54 ;
   RECT 23.18 639.54 933.28 641.25 ;
   RECT 23.18 641.25 933.28 642.96 ;
   RECT 23.18 642.96 933.28 644.67 ;
   RECT 23.18 644.67 933.28 646.38 ;
   RECT 23.18 646.38 933.28 648.09 ;
   RECT 23.18 648.09 933.28 649.8 ;
   RECT 23.18 649.8 933.28 651.51 ;
   RECT 23.18 651.51 933.28 653.22 ;
   RECT 23.18 653.22 933.28 654.93 ;
   RECT 23.18 654.93 933.28 656.64 ;
   RECT 23.18 656.64 933.28 658.35 ;
   RECT 23.18 658.35 933.28 660.06 ;
   RECT 23.18 660.06 933.28 661.77 ;
   RECT 23.18 661.77 933.28 663.48 ;
   RECT 23.18 663.48 933.28 665.19 ;
   RECT 23.18 665.19 933.28 666.9 ;
   RECT 23.18 666.9 933.28 668.61 ;
   RECT 23.18 668.61 933.28 670.32 ;
   RECT 23.18 670.32 933.28 672.03 ;
   RECT 23.18 672.03 933.28 673.74 ;
   RECT 23.18 673.74 933.28 675.45 ;
   RECT 23.18 675.45 933.28 677.16 ;
   RECT 23.18 677.16 933.28 678.87 ;
   RECT 23.18 678.87 933.28 680.58 ;
   RECT 23.18 680.58 933.28 682.29 ;
   RECT 23.18 682.29 933.28 684.0 ;
   RECT 23.18 684.0 933.28 685.71 ;
   RECT 23.18 685.71 933.28 687.42 ;
   RECT 23.18 687.42 933.28 689.13 ;
   RECT 23.18 689.13 933.28 690.84 ;
   RECT 23.18 690.84 933.28 692.55 ;
   RECT 23.18 692.55 933.28 694.26 ;
   RECT 23.18 694.26 933.28 695.97 ;
   RECT 23.18 695.97 933.28 697.68 ;
   RECT 23.18 697.68 933.28 699.39 ;
   RECT 23.18 699.39 933.28 701.1 ;
   RECT 23.18 701.1 933.28 702.81 ;
   RECT 23.18 702.81 933.28 704.52 ;
   RECT 23.18 704.52 933.28 706.23 ;
   RECT 23.18 706.23 933.28 707.94 ;
   RECT 23.18 707.94 933.28 709.65 ;
   RECT 23.18 709.65 933.28 711.36 ;
   RECT 23.18 711.36 933.28 713.07 ;
   RECT 23.18 713.07 933.28 714.78 ;
   RECT 23.18 714.78 933.28 716.49 ;
   RECT 23.18 716.49 933.28 718.2 ;
   RECT 23.18 718.2 933.28 719.91 ;
   RECT 23.18 719.91 933.28 721.62 ;
   RECT 23.18 721.62 933.28 723.33 ;
   RECT 23.18 723.33 933.28 725.04 ;
   RECT 23.18 725.04 933.28 726.75 ;
   RECT 23.18 726.75 933.28 728.46 ;
   RECT 23.18 728.46 933.28 730.17 ;
   RECT 23.18 730.17 933.28 731.88 ;
   RECT 23.18 731.88 933.28 733.59 ;
   RECT 23.18 733.59 933.28 735.3 ;
   RECT 23.18 735.3 933.28 737.01 ;
   RECT 23.18 737.01 933.28 738.72 ;
   RECT 23.18 738.72 933.28 740.43 ;
   RECT 23.18 740.43 933.28 742.14 ;
   RECT 23.18 742.14 933.28 743.85 ;
   RECT 23.18 743.85 933.28 745.56 ;
   RECT 23.18 745.56 933.28 747.27 ;
   RECT 23.18 747.27 933.28 748.98 ;
   RECT 23.18 748.98 933.28 750.69 ;
   RECT 23.18 750.69 933.28 752.4 ;
   RECT 23.18 752.4 933.28 754.11 ;
   RECT 23.18 754.11 933.28 755.82 ;
   RECT 23.18 755.82 933.28 757.53 ;
   RECT 23.18 757.53 933.28 759.24 ;
   RECT 23.18 759.24 933.28 760.95 ;
   RECT 23.18 760.95 933.28 762.66 ;
   RECT 23.18 762.66 933.28 764.37 ;
   RECT 23.18 764.37 933.28 766.08 ;
   RECT 23.18 766.08 933.28 767.79 ;
   RECT 23.18 767.79 933.28 769.5 ;
   RECT 23.18 769.5 933.28 771.21 ;
   RECT 23.18 771.21 933.28 772.92 ;
   RECT 23.18 772.92 933.28 774.63 ;
   RECT 23.18 774.63 933.28 776.34 ;
   RECT 23.18 776.34 933.28 778.05 ;
   RECT 23.18 778.05 933.28 779.76 ;
   RECT 23.18 779.76 933.28 781.47 ;
   RECT 23.18 781.47 933.28 783.18 ;
   RECT 23.18 783.18 933.28 784.89 ;
   RECT 23.18 784.89 933.28 786.6 ;
   RECT 23.18 786.6 933.28 788.31 ;
   RECT 23.18 788.31 933.28 790.02 ;
   RECT 23.18 790.02 933.28 791.73 ;
   RECT 23.18 791.73 933.28 793.44 ;
   RECT 23.18 793.44 933.28 795.15 ;
   RECT 23.18 795.15 933.28 796.86 ;
   RECT 23.18 796.86 933.28 798.57 ;
   RECT 23.18 798.57 933.28 800.28 ;
   RECT 23.18 800.28 933.28 801.99 ;
   RECT 23.18 801.99 933.28 803.7 ;
   RECT 23.18 803.7 933.28 805.41 ;
   RECT 23.18 805.41 933.28 807.12 ;
   RECT 23.18 807.12 933.28 808.83 ;
   RECT 23.18 808.83 933.28 810.54 ;
   RECT 23.18 810.54 933.28 812.25 ;
   RECT 23.18 812.25 933.28 813.96 ;
   RECT 23.18 813.96 933.28 815.67 ;
   RECT 23.18 815.67 933.28 817.38 ;
   RECT 23.18 817.38 933.28 819.09 ;
   RECT 23.18 819.09 933.28 820.8 ;
   RECT 23.18 820.8 933.28 822.51 ;
   RECT 23.18 822.51 933.28 824.22 ;
   RECT 23.18 824.22 933.28 825.93 ;
   RECT 23.18 825.93 933.28 827.64 ;
   RECT 23.18 827.64 933.28 829.35 ;
   RECT 23.18 829.35 933.28 831.06 ;
   RECT 23.18 831.06 933.28 832.77 ;
   RECT 23.18 832.77 933.28 834.48 ;
   RECT 23.18 834.48 933.28 836.19 ;
   RECT 23.18 836.19 933.28 837.9 ;
   RECT 23.18 837.9 933.28 839.61 ;
   RECT 23.18 839.61 933.28 841.32 ;
   RECT 23.18 841.32 933.28 843.03 ;
   RECT 23.18 843.03 933.28 844.74 ;
   RECT 23.18 844.74 933.28 846.45 ;
   RECT 23.18 846.45 933.28 848.16 ;
   RECT 23.18 848.16 933.28 849.87 ;
   RECT 23.18 849.87 933.28 851.58 ;
   RECT 23.18 851.58 933.28 853.29 ;
   RECT 23.18 853.29 933.28 855.0 ;
   RECT 23.18 855.0 933.28 856.71 ;
   RECT 23.18 856.71 933.28 858.42 ;
   RECT 23.18 858.42 933.28 860.13 ;
   RECT 23.18 860.13 933.28 861.84 ;
   RECT 23.18 861.84 933.28 863.55 ;
   RECT 23.18 863.55 933.28 865.26 ;
   RECT 23.18 865.26 933.28 866.97 ;
   RECT 23.18 866.97 933.28 868.68 ;
   RECT 23.18 868.68 933.28 870.39 ;
   RECT 23.18 870.39 933.28 872.1 ;
   RECT 23.18 872.1 933.28 873.81 ;
   RECT 23.18 873.81 933.28 875.52 ;
   RECT 23.18 875.52 933.28 877.23 ;
   RECT 23.18 877.23 933.28 878.94 ;
  LAYER via2 ;
   RECT 23.18 0.0 933.28 1.71 ;
   RECT 23.18 1.71 933.28 3.42 ;
   RECT 23.18 3.42 933.28 5.13 ;
   RECT 23.18 5.13 933.28 6.84 ;
   RECT 23.18 6.84 933.28 8.55 ;
   RECT 23.18 8.55 933.28 10.26 ;
   RECT 23.18 10.26 933.28 11.97 ;
   RECT 23.18 11.97 933.28 13.68 ;
   RECT 23.18 13.68 933.28 15.39 ;
   RECT 23.18 15.39 933.28 17.1 ;
   RECT 23.18 17.1 933.28 18.81 ;
   RECT 23.18 18.81 933.28 20.52 ;
   RECT 23.18 20.52 933.28 22.23 ;
   RECT 23.18 22.23 933.28 23.94 ;
   RECT 23.18 23.94 933.28 25.65 ;
   RECT 23.18 25.65 933.28 27.36 ;
   RECT 23.18 27.36 933.28 29.07 ;
   RECT 23.18 29.07 933.28 30.78 ;
   RECT 23.18 30.78 933.28 32.49 ;
   RECT 23.18 32.49 933.28 34.2 ;
   RECT 23.18 34.2 933.28 35.91 ;
   RECT 23.18 35.91 933.28 37.62 ;
   RECT 23.18 37.62 933.28 39.33 ;
   RECT 23.18 39.33 933.28 41.04 ;
   RECT 23.18 41.04 933.28 42.75 ;
   RECT 23.18 42.75 933.28 44.46 ;
   RECT 23.18 44.46 933.28 46.17 ;
   RECT 23.18 46.17 933.28 47.88 ;
   RECT 23.18 47.88 933.28 49.59 ;
   RECT 23.18 49.59 933.28 51.3 ;
   RECT 23.18 51.3 933.28 53.01 ;
   RECT 23.18 53.01 933.28 54.72 ;
   RECT 23.18 54.72 933.28 56.43 ;
   RECT 23.18 56.43 933.28 58.14 ;
   RECT 23.18 58.14 933.28 59.85 ;
   RECT 23.18 59.85 933.28 61.56 ;
   RECT 23.18 61.56 933.28 63.27 ;
   RECT 23.18 63.27 933.28 64.98 ;
   RECT 23.18 64.98 933.28 66.69 ;
   RECT 23.18 66.69 933.28 68.4 ;
   RECT 23.18 68.4 933.28 70.11 ;
   RECT 23.18 70.11 933.28 71.82 ;
   RECT 23.18 71.82 933.28 73.53 ;
   RECT 23.18 73.53 933.28 75.24 ;
   RECT 23.18 75.24 933.28 76.95 ;
   RECT 23.18 76.95 933.28 78.66 ;
   RECT 23.18 78.66 933.28 80.37 ;
   RECT 23.18 80.37 933.28 82.08 ;
   RECT 23.18 82.08 933.28 83.79 ;
   RECT 23.18 83.79 933.28 85.5 ;
   RECT 23.18 85.5 933.28 87.21 ;
   RECT 23.18 87.21 933.28 88.92 ;
   RECT 23.18 88.92 933.28 90.63 ;
   RECT 23.18 90.63 933.28 92.34 ;
   RECT 23.18 92.34 933.28 94.05 ;
   RECT 23.18 94.05 933.28 95.76 ;
   RECT 23.18 95.76 933.28 97.47 ;
   RECT 23.18 97.47 933.28 99.18 ;
   RECT 23.18 99.18 933.28 100.89 ;
   RECT 23.18 100.89 933.28 102.6 ;
   RECT 23.18 102.6 933.28 104.31 ;
   RECT 23.18 104.31 933.28 106.02 ;
   RECT 23.18 106.02 933.28 107.73 ;
   RECT 23.18 107.73 933.28 109.44 ;
   RECT 23.18 109.44 933.28 111.15 ;
   RECT 23.18 111.15 933.28 112.86 ;
   RECT 23.18 112.86 933.28 114.57 ;
   RECT 23.18 114.57 933.28 116.28 ;
   RECT 23.18 116.28 933.28 117.99 ;
   RECT 23.18 117.99 933.28 119.7 ;
   RECT 23.18 119.7 933.28 121.41 ;
   RECT 23.18 121.41 933.28 123.12 ;
   RECT 23.18 123.12 933.28 124.83 ;
   RECT 23.18 124.83 933.28 126.54 ;
   RECT 23.18 126.54 933.28 128.25 ;
   RECT 23.18 128.25 933.28 129.96 ;
   RECT 23.18 129.96 933.28 131.67 ;
   RECT 23.18 131.67 933.28 133.38 ;
   RECT 23.18 133.38 933.28 135.09 ;
   RECT 23.18 135.09 933.28 136.8 ;
   RECT 23.18 136.8 933.28 138.51 ;
   RECT 23.18 138.51 933.28 140.22 ;
   RECT 23.18 140.22 933.28 141.93 ;
   RECT 23.18 141.93 933.28 143.64 ;
   RECT 23.18 143.64 933.28 145.35 ;
   RECT 23.18 145.35 933.28 147.06 ;
   RECT 23.18 147.06 933.28 148.77 ;
   RECT 23.18 148.77 933.28 150.48 ;
   RECT 23.18 150.48 933.28 152.19 ;
   RECT 23.18 152.19 933.28 153.9 ;
   RECT 23.18 153.9 933.28 155.61 ;
   RECT 23.18 155.61 933.28 157.32 ;
   RECT 23.18 157.32 933.28 159.03 ;
   RECT 23.18 159.03 933.28 160.74 ;
   RECT 23.18 160.74 933.28 162.45 ;
   RECT 23.18 162.45 933.28 164.16 ;
   RECT 23.18 164.16 933.28 165.87 ;
   RECT 23.18 165.87 933.28 167.58 ;
   RECT 23.18 167.58 933.28 169.29 ;
   RECT 23.18 169.29 933.28 171.0 ;
   RECT 23.18 171.0 933.28 172.71 ;
   RECT 23.18 172.71 933.28 174.42 ;
   RECT 23.18 174.42 933.28 176.13 ;
   RECT 23.18 176.13 933.28 177.84 ;
   RECT 23.18 177.84 933.28 179.55 ;
   RECT 23.18 179.55 933.28 181.26 ;
   RECT 23.18 181.26 933.28 182.97 ;
   RECT 23.18 182.97 933.28 184.68 ;
   RECT 23.18 184.68 933.28 186.39 ;
   RECT 23.18 186.39 933.28 188.1 ;
   RECT 23.18 188.1 933.28 189.81 ;
   RECT 23.18 189.81 933.28 191.52 ;
   RECT 23.18 191.52 933.28 193.23 ;
   RECT 23.18 193.23 933.28 194.94 ;
   RECT 23.18 194.94 933.28 196.65 ;
   RECT 23.18 196.65 933.28 198.36 ;
   RECT 23.18 198.36 933.28 200.07 ;
   RECT 23.18 200.07 933.28 201.78 ;
   RECT 23.18 201.78 933.28 203.49 ;
   RECT 23.18 203.49 933.28 205.2 ;
   RECT 23.18 205.2 933.28 206.91 ;
   RECT 23.18 206.91 933.28 208.62 ;
   RECT 23.18 208.62 933.28 210.33 ;
   RECT 23.18 210.33 933.28 212.04 ;
   RECT 23.18 212.04 933.28 213.75 ;
   RECT 23.18 213.75 933.28 215.46 ;
   RECT 23.18 215.46 933.28 217.17 ;
   RECT 23.18 217.17 933.28 218.88 ;
   RECT 23.18 218.88 933.28 220.59 ;
   RECT 23.18 220.59 933.28 222.3 ;
   RECT 23.18 222.3 933.28 224.01 ;
   RECT 23.18 224.01 933.28 225.72 ;
   RECT 23.18 225.72 933.28 227.43 ;
   RECT 23.18 227.43 933.28 229.14 ;
   RECT 23.18 229.14 933.28 230.85 ;
   RECT 23.18 230.85 933.28 232.56 ;
   RECT 23.18 232.56 933.28 234.27 ;
   RECT 23.18 234.27 933.28 235.98 ;
   RECT 23.18 235.98 933.28 237.69 ;
   RECT 23.18 237.69 933.28 239.4 ;
   RECT 23.18 239.4 933.28 241.11 ;
   RECT 23.18 241.11 933.28 242.82 ;
   RECT 23.18 242.82 933.28 244.53 ;
   RECT 23.18 244.53 933.28 246.24 ;
   RECT 23.18 246.24 933.28 247.95 ;
   RECT 23.18 247.95 933.28 249.66 ;
   RECT 23.18 249.66 933.28 251.37 ;
   RECT 23.18 251.37 933.28 253.08 ;
   RECT 23.18 253.08 933.28 254.79 ;
   RECT 23.18 254.79 933.28 256.5 ;
   RECT 23.18 256.5 933.28 258.21 ;
   RECT 23.18 258.21 933.28 259.92 ;
   RECT 23.18 259.92 933.28 261.63 ;
   RECT 23.18 261.63 933.28 263.34 ;
   RECT 23.18 263.34 933.28 265.05 ;
   RECT 23.18 265.05 933.28 266.76 ;
   RECT 23.18 266.76 933.28 268.47 ;
   RECT 23.18 268.47 933.28 270.18 ;
   RECT 23.18 270.18 933.28 271.89 ;
   RECT 23.18 271.89 933.28 273.6 ;
   RECT 23.18 273.6 933.28 275.31 ;
   RECT 23.18 275.31 933.28 277.02 ;
   RECT 23.18 277.02 933.28 278.73 ;
   RECT 23.18 278.73 933.28 280.44 ;
   RECT 23.18 280.44 933.28 282.15 ;
   RECT 23.18 282.15 933.28 283.86 ;
   RECT 23.18 283.86 933.28 285.57 ;
   RECT 23.18 285.57 933.28 287.28 ;
   RECT 23.18 287.28 933.28 288.99 ;
   RECT 23.18 288.99 933.28 290.7 ;
   RECT 23.18 290.7 933.28 292.41 ;
   RECT 23.18 292.41 933.28 294.12 ;
   RECT 23.18 294.12 933.28 295.83 ;
   RECT 23.18 295.83 933.28 297.54 ;
   RECT 23.18 297.54 933.28 299.25 ;
   RECT 23.18 299.25 933.28 300.96 ;
   RECT 23.18 300.96 933.28 302.67 ;
   RECT 23.18 302.67 933.28 304.38 ;
   RECT 23.18 304.38 933.28 306.09 ;
   RECT 23.18 306.09 933.28 307.8 ;
   RECT 23.18 307.8 933.28 309.51 ;
   RECT 23.18 309.51 933.28 311.22 ;
   RECT 23.18 311.22 933.28 312.93 ;
   RECT 23.18 312.93 933.28 314.64 ;
   RECT 23.18 314.64 933.28 316.35 ;
   RECT 23.18 316.35 933.28 318.06 ;
   RECT 23.18 318.06 933.28 319.77 ;
   RECT 23.18 319.77 933.28 321.48 ;
   RECT 23.18 321.48 933.28 323.19 ;
   RECT 23.18 323.19 933.28 324.9 ;
   RECT 23.18 324.9 933.28 326.61 ;
   RECT 23.18 326.61 933.28 328.32 ;
   RECT 23.18 328.32 933.28 330.03 ;
   RECT 23.18 330.03 933.28 331.74 ;
   RECT 23.18 331.74 933.28 333.45 ;
   RECT 23.18 333.45 933.28 335.16 ;
   RECT 23.18 335.16 933.28 336.87 ;
   RECT 23.18 336.87 933.28 338.58 ;
   RECT 23.18 338.58 933.28 340.29 ;
   RECT 23.18 340.29 933.28 342.0 ;
   RECT 23.18 342.0 933.28 343.71 ;
   RECT 23.18 343.71 933.28 345.42 ;
   RECT 23.18 345.42 933.28 347.13 ;
   RECT 23.18 347.13 933.28 348.84 ;
   RECT 23.18 348.84 933.28 350.55 ;
   RECT 23.18 350.55 933.28 352.26 ;
   RECT 23.18 352.26 933.28 353.97 ;
   RECT 23.18 353.97 933.28 355.68 ;
   RECT 23.18 355.68 933.28 357.39 ;
   RECT 23.18 357.39 933.28 359.1 ;
   RECT 23.18 359.1 933.28 360.81 ;
   RECT 23.18 360.81 933.28 362.52 ;
   RECT 23.18 362.52 933.28 364.23 ;
   RECT 23.18 364.23 933.28 365.94 ;
   RECT 23.18 365.94 933.28 367.65 ;
   RECT 23.18 367.65 933.28 369.36 ;
   RECT 23.18 369.36 933.28 371.07 ;
   RECT 23.18 371.07 933.28 372.78 ;
   RECT 23.18 372.78 933.28 374.49 ;
   RECT 23.18 374.49 933.28 376.2 ;
   RECT 23.18 376.2 933.28 377.91 ;
   RECT 23.18 377.91 933.28 379.62 ;
   RECT 23.18 379.62 933.28 381.33 ;
   RECT 23.18 381.33 933.28 383.04 ;
   RECT 23.18 383.04 933.28 384.75 ;
   RECT 23.18 384.75 933.28 386.46 ;
   RECT 23.18 386.46 933.28 388.17 ;
   RECT 23.18 388.17 933.28 389.88 ;
   RECT 23.18 389.88 933.28 391.59 ;
   RECT 23.18 391.59 933.28 393.3 ;
   RECT 23.18 393.3 933.28 395.01 ;
   RECT 23.18 395.01 933.28 396.72 ;
   RECT 23.18 396.72 933.28 398.43 ;
   RECT 23.18 398.43 933.28 400.14 ;
   RECT 23.18 400.14 933.28 401.85 ;
   RECT 23.18 401.85 933.28 403.56 ;
   RECT 23.18 403.56 933.28 405.27 ;
   RECT 23.18 405.27 933.28 406.98 ;
   RECT 23.18 406.98 933.28 408.69 ;
   RECT 23.18 408.69 933.28 410.4 ;
   RECT 23.18 410.4 933.28 412.11 ;
   RECT 23.18 412.11 933.28 413.82 ;
   RECT 23.18 413.82 933.28 415.53 ;
   RECT 23.18 415.53 933.28 417.24 ;
   RECT 23.18 417.24 933.28 418.95 ;
   RECT 23.18 418.95 933.28 420.66 ;
   RECT 23.18 420.66 933.28 422.37 ;
   RECT 23.18 422.37 933.28 424.08 ;
   RECT 23.18 424.08 933.28 425.79 ;
   RECT 23.18 425.79 933.28 427.5 ;
   RECT 23.18 427.5 933.28 429.21 ;
   RECT 23.18 429.21 933.28 430.92 ;
   RECT 0.0 430.92 933.28 432.63 ;
   RECT 0.0 432.63 933.28 434.34 ;
   RECT 0.0 434.34 933.28 436.05 ;
   RECT 0.0 436.05 933.28 437.76 ;
   RECT 0.0 437.76 933.28 439.47 ;
   RECT 0.0 439.47 933.28 441.18 ;
   RECT 0.0 441.18 933.28 442.89 ;
   RECT 0.0 442.89 933.28 444.6 ;
   RECT 0.0 444.6 933.28 446.31 ;
   RECT 0.0 446.31 933.28 448.02 ;
   RECT 0.0 448.02 933.28 449.73 ;
   RECT 0.0 449.73 933.28 451.44 ;
   RECT 0.0 451.44 933.28 453.15 ;
   RECT 0.0 453.15 933.28 454.86 ;
   RECT 0.0 454.86 933.28 456.57 ;
   RECT 0.0 456.57 933.28 458.28 ;
   RECT 0.0 458.28 933.28 459.99 ;
   RECT 23.18 459.99 933.28 461.7 ;
   RECT 23.18 461.7 933.28 463.41 ;
   RECT 23.18 463.41 933.28 465.12 ;
   RECT 23.18 465.12 933.28 466.83 ;
   RECT 23.18 466.83 933.28 468.54 ;
   RECT 23.18 468.54 933.28 470.25 ;
   RECT 23.18 470.25 933.28 471.96 ;
   RECT 23.18 471.96 933.28 473.67 ;
   RECT 23.18 473.67 933.28 475.38 ;
   RECT 23.18 475.38 933.28 477.09 ;
   RECT 23.18 477.09 933.28 478.8 ;
   RECT 23.18 478.8 933.28 480.51 ;
   RECT 23.18 480.51 933.28 482.22 ;
   RECT 23.18 482.22 933.28 483.93 ;
   RECT 23.18 483.93 933.28 485.64 ;
   RECT 23.18 485.64 933.28 487.35 ;
   RECT 23.18 487.35 933.28 489.06 ;
   RECT 23.18 489.06 933.28 490.77 ;
   RECT 23.18 490.77 933.28 492.48 ;
   RECT 23.18 492.48 933.28 494.19 ;
   RECT 23.18 494.19 933.28 495.9 ;
   RECT 23.18 495.9 933.28 497.61 ;
   RECT 23.18 497.61 933.28 499.32 ;
   RECT 23.18 499.32 933.28 501.03 ;
   RECT 23.18 501.03 933.28 502.74 ;
   RECT 23.18 502.74 933.28 504.45 ;
   RECT 23.18 504.45 933.28 506.16 ;
   RECT 23.18 506.16 933.28 507.87 ;
   RECT 23.18 507.87 933.28 509.58 ;
   RECT 23.18 509.58 933.28 511.29 ;
   RECT 23.18 511.29 933.28 513.0 ;
   RECT 23.18 513.0 933.28 514.71 ;
   RECT 23.18 514.71 933.28 516.42 ;
   RECT 23.18 516.42 933.28 518.13 ;
   RECT 23.18 518.13 933.28 519.84 ;
   RECT 23.18 519.84 933.28 521.55 ;
   RECT 23.18 521.55 933.28 523.26 ;
   RECT 23.18 523.26 933.28 524.97 ;
   RECT 23.18 524.97 933.28 526.68 ;
   RECT 23.18 526.68 933.28 528.39 ;
   RECT 23.18 528.39 933.28 530.1 ;
   RECT 23.18 530.1 933.28 531.81 ;
   RECT 23.18 531.81 933.28 533.52 ;
   RECT 23.18 533.52 933.28 535.23 ;
   RECT 23.18 535.23 933.28 536.94 ;
   RECT 23.18 536.94 933.28 538.65 ;
   RECT 23.18 538.65 933.28 540.36 ;
   RECT 23.18 540.36 933.28 542.07 ;
   RECT 23.18 542.07 933.28 543.78 ;
   RECT 23.18 543.78 933.28 545.49 ;
   RECT 23.18 545.49 933.28 547.2 ;
   RECT 23.18 547.2 933.28 548.91 ;
   RECT 23.18 548.91 933.28 550.62 ;
   RECT 23.18 550.62 933.28 552.33 ;
   RECT 23.18 552.33 933.28 554.04 ;
   RECT 23.18 554.04 933.28 555.75 ;
   RECT 23.18 555.75 933.28 557.46 ;
   RECT 23.18 557.46 933.28 559.17 ;
   RECT 23.18 559.17 933.28 560.88 ;
   RECT 23.18 560.88 933.28 562.59 ;
   RECT 23.18 562.59 933.28 564.3 ;
   RECT 23.18 564.3 933.28 566.01 ;
   RECT 23.18 566.01 933.28 567.72 ;
   RECT 23.18 567.72 933.28 569.43 ;
   RECT 23.18 569.43 933.28 571.14 ;
   RECT 23.18 571.14 933.28 572.85 ;
   RECT 23.18 572.85 933.28 574.56 ;
   RECT 23.18 574.56 933.28 576.27 ;
   RECT 23.18 576.27 933.28 577.98 ;
   RECT 23.18 577.98 933.28 579.69 ;
   RECT 23.18 579.69 933.28 581.4 ;
   RECT 23.18 581.4 933.28 583.11 ;
   RECT 23.18 583.11 933.28 584.82 ;
   RECT 23.18 584.82 933.28 586.53 ;
   RECT 23.18 586.53 933.28 588.24 ;
   RECT 23.18 588.24 933.28 589.95 ;
   RECT 23.18 589.95 933.28 591.66 ;
   RECT 23.18 591.66 933.28 593.37 ;
   RECT 23.18 593.37 933.28 595.08 ;
   RECT 23.18 595.08 933.28 596.79 ;
   RECT 23.18 596.79 933.28 598.5 ;
   RECT 23.18 598.5 933.28 600.21 ;
   RECT 23.18 600.21 933.28 601.92 ;
   RECT 23.18 601.92 933.28 603.63 ;
   RECT 23.18 603.63 933.28 605.34 ;
   RECT 23.18 605.34 933.28 607.05 ;
   RECT 23.18 607.05 933.28 608.76 ;
   RECT 23.18 608.76 933.28 610.47 ;
   RECT 23.18 610.47 933.28 612.18 ;
   RECT 23.18 612.18 933.28 613.89 ;
   RECT 23.18 613.89 933.28 615.6 ;
   RECT 23.18 615.6 933.28 617.31 ;
   RECT 23.18 617.31 933.28 619.02 ;
   RECT 23.18 619.02 933.28 620.73 ;
   RECT 23.18 620.73 933.28 622.44 ;
   RECT 23.18 622.44 933.28 624.15 ;
   RECT 23.18 624.15 933.28 625.86 ;
   RECT 23.18 625.86 933.28 627.57 ;
   RECT 23.18 627.57 933.28 629.28 ;
   RECT 23.18 629.28 933.28 630.99 ;
   RECT 23.18 630.99 933.28 632.7 ;
   RECT 23.18 632.7 933.28 634.41 ;
   RECT 23.18 634.41 933.28 636.12 ;
   RECT 23.18 636.12 933.28 637.83 ;
   RECT 23.18 637.83 933.28 639.54 ;
   RECT 23.18 639.54 933.28 641.25 ;
   RECT 23.18 641.25 933.28 642.96 ;
   RECT 23.18 642.96 933.28 644.67 ;
   RECT 23.18 644.67 933.28 646.38 ;
   RECT 23.18 646.38 933.28 648.09 ;
   RECT 23.18 648.09 933.28 649.8 ;
   RECT 23.18 649.8 933.28 651.51 ;
   RECT 23.18 651.51 933.28 653.22 ;
   RECT 23.18 653.22 933.28 654.93 ;
   RECT 23.18 654.93 933.28 656.64 ;
   RECT 23.18 656.64 933.28 658.35 ;
   RECT 23.18 658.35 933.28 660.06 ;
   RECT 23.18 660.06 933.28 661.77 ;
   RECT 23.18 661.77 933.28 663.48 ;
   RECT 23.18 663.48 933.28 665.19 ;
   RECT 23.18 665.19 933.28 666.9 ;
   RECT 23.18 666.9 933.28 668.61 ;
   RECT 23.18 668.61 933.28 670.32 ;
   RECT 23.18 670.32 933.28 672.03 ;
   RECT 23.18 672.03 933.28 673.74 ;
   RECT 23.18 673.74 933.28 675.45 ;
   RECT 23.18 675.45 933.28 677.16 ;
   RECT 23.18 677.16 933.28 678.87 ;
   RECT 23.18 678.87 933.28 680.58 ;
   RECT 23.18 680.58 933.28 682.29 ;
   RECT 23.18 682.29 933.28 684.0 ;
   RECT 23.18 684.0 933.28 685.71 ;
   RECT 23.18 685.71 933.28 687.42 ;
   RECT 23.18 687.42 933.28 689.13 ;
   RECT 23.18 689.13 933.28 690.84 ;
   RECT 23.18 690.84 933.28 692.55 ;
   RECT 23.18 692.55 933.28 694.26 ;
   RECT 23.18 694.26 933.28 695.97 ;
   RECT 23.18 695.97 933.28 697.68 ;
   RECT 23.18 697.68 933.28 699.39 ;
   RECT 23.18 699.39 933.28 701.1 ;
   RECT 23.18 701.1 933.28 702.81 ;
   RECT 23.18 702.81 933.28 704.52 ;
   RECT 23.18 704.52 933.28 706.23 ;
   RECT 23.18 706.23 933.28 707.94 ;
   RECT 23.18 707.94 933.28 709.65 ;
   RECT 23.18 709.65 933.28 711.36 ;
   RECT 23.18 711.36 933.28 713.07 ;
   RECT 23.18 713.07 933.28 714.78 ;
   RECT 23.18 714.78 933.28 716.49 ;
   RECT 23.18 716.49 933.28 718.2 ;
   RECT 23.18 718.2 933.28 719.91 ;
   RECT 23.18 719.91 933.28 721.62 ;
   RECT 23.18 721.62 933.28 723.33 ;
   RECT 23.18 723.33 933.28 725.04 ;
   RECT 23.18 725.04 933.28 726.75 ;
   RECT 23.18 726.75 933.28 728.46 ;
   RECT 23.18 728.46 933.28 730.17 ;
   RECT 23.18 730.17 933.28 731.88 ;
   RECT 23.18 731.88 933.28 733.59 ;
   RECT 23.18 733.59 933.28 735.3 ;
   RECT 23.18 735.3 933.28 737.01 ;
   RECT 23.18 737.01 933.28 738.72 ;
   RECT 23.18 738.72 933.28 740.43 ;
   RECT 23.18 740.43 933.28 742.14 ;
   RECT 23.18 742.14 933.28 743.85 ;
   RECT 23.18 743.85 933.28 745.56 ;
   RECT 23.18 745.56 933.28 747.27 ;
   RECT 23.18 747.27 933.28 748.98 ;
   RECT 23.18 748.98 933.28 750.69 ;
   RECT 23.18 750.69 933.28 752.4 ;
   RECT 23.18 752.4 933.28 754.11 ;
   RECT 23.18 754.11 933.28 755.82 ;
   RECT 23.18 755.82 933.28 757.53 ;
   RECT 23.18 757.53 933.28 759.24 ;
   RECT 23.18 759.24 933.28 760.95 ;
   RECT 23.18 760.95 933.28 762.66 ;
   RECT 23.18 762.66 933.28 764.37 ;
   RECT 23.18 764.37 933.28 766.08 ;
   RECT 23.18 766.08 933.28 767.79 ;
   RECT 23.18 767.79 933.28 769.5 ;
   RECT 23.18 769.5 933.28 771.21 ;
   RECT 23.18 771.21 933.28 772.92 ;
   RECT 23.18 772.92 933.28 774.63 ;
   RECT 23.18 774.63 933.28 776.34 ;
   RECT 23.18 776.34 933.28 778.05 ;
   RECT 23.18 778.05 933.28 779.76 ;
   RECT 23.18 779.76 933.28 781.47 ;
   RECT 23.18 781.47 933.28 783.18 ;
   RECT 23.18 783.18 933.28 784.89 ;
   RECT 23.18 784.89 933.28 786.6 ;
   RECT 23.18 786.6 933.28 788.31 ;
   RECT 23.18 788.31 933.28 790.02 ;
   RECT 23.18 790.02 933.28 791.73 ;
   RECT 23.18 791.73 933.28 793.44 ;
   RECT 23.18 793.44 933.28 795.15 ;
   RECT 23.18 795.15 933.28 796.86 ;
   RECT 23.18 796.86 933.28 798.57 ;
   RECT 23.18 798.57 933.28 800.28 ;
   RECT 23.18 800.28 933.28 801.99 ;
   RECT 23.18 801.99 933.28 803.7 ;
   RECT 23.18 803.7 933.28 805.41 ;
   RECT 23.18 805.41 933.28 807.12 ;
   RECT 23.18 807.12 933.28 808.83 ;
   RECT 23.18 808.83 933.28 810.54 ;
   RECT 23.18 810.54 933.28 812.25 ;
   RECT 23.18 812.25 933.28 813.96 ;
   RECT 23.18 813.96 933.28 815.67 ;
   RECT 23.18 815.67 933.28 817.38 ;
   RECT 23.18 817.38 933.28 819.09 ;
   RECT 23.18 819.09 933.28 820.8 ;
   RECT 23.18 820.8 933.28 822.51 ;
   RECT 23.18 822.51 933.28 824.22 ;
   RECT 23.18 824.22 933.28 825.93 ;
   RECT 23.18 825.93 933.28 827.64 ;
   RECT 23.18 827.64 933.28 829.35 ;
   RECT 23.18 829.35 933.28 831.06 ;
   RECT 23.18 831.06 933.28 832.77 ;
   RECT 23.18 832.77 933.28 834.48 ;
   RECT 23.18 834.48 933.28 836.19 ;
   RECT 23.18 836.19 933.28 837.9 ;
   RECT 23.18 837.9 933.28 839.61 ;
   RECT 23.18 839.61 933.28 841.32 ;
   RECT 23.18 841.32 933.28 843.03 ;
   RECT 23.18 843.03 933.28 844.74 ;
   RECT 23.18 844.74 933.28 846.45 ;
   RECT 23.18 846.45 933.28 848.16 ;
   RECT 23.18 848.16 933.28 849.87 ;
   RECT 23.18 849.87 933.28 851.58 ;
   RECT 23.18 851.58 933.28 853.29 ;
   RECT 23.18 853.29 933.28 855.0 ;
   RECT 23.18 855.0 933.28 856.71 ;
   RECT 23.18 856.71 933.28 858.42 ;
   RECT 23.18 858.42 933.28 860.13 ;
   RECT 23.18 860.13 933.28 861.84 ;
   RECT 23.18 861.84 933.28 863.55 ;
   RECT 23.18 863.55 933.28 865.26 ;
   RECT 23.18 865.26 933.28 866.97 ;
   RECT 23.18 866.97 933.28 868.68 ;
   RECT 23.18 868.68 933.28 870.39 ;
   RECT 23.18 870.39 933.28 872.1 ;
   RECT 23.18 872.1 933.28 873.81 ;
   RECT 23.18 873.81 933.28 875.52 ;
   RECT 23.18 875.52 933.28 877.23 ;
   RECT 23.18 877.23 933.28 878.94 ;
  LAYER metal3 ;
   RECT 23.18 0.0 933.28 1.71 ;
   RECT 23.18 1.71 933.28 3.42 ;
   RECT 23.18 3.42 933.28 5.13 ;
   RECT 23.18 5.13 933.28 6.84 ;
   RECT 23.18 6.84 933.28 8.55 ;
   RECT 23.18 8.55 933.28 10.26 ;
   RECT 23.18 10.26 933.28 11.97 ;
   RECT 23.18 11.97 933.28 13.68 ;
   RECT 23.18 13.68 933.28 15.39 ;
   RECT 23.18 15.39 933.28 17.1 ;
   RECT 23.18 17.1 933.28 18.81 ;
   RECT 23.18 18.81 933.28 20.52 ;
   RECT 23.18 20.52 933.28 22.23 ;
   RECT 23.18 22.23 933.28 23.94 ;
   RECT 23.18 23.94 933.28 25.65 ;
   RECT 23.18 25.65 933.28 27.36 ;
   RECT 23.18 27.36 933.28 29.07 ;
   RECT 23.18 29.07 933.28 30.78 ;
   RECT 23.18 30.78 933.28 32.49 ;
   RECT 23.18 32.49 933.28 34.2 ;
   RECT 23.18 34.2 933.28 35.91 ;
   RECT 23.18 35.91 933.28 37.62 ;
   RECT 23.18 37.62 933.28 39.33 ;
   RECT 23.18 39.33 933.28 41.04 ;
   RECT 23.18 41.04 933.28 42.75 ;
   RECT 23.18 42.75 933.28 44.46 ;
   RECT 23.18 44.46 933.28 46.17 ;
   RECT 23.18 46.17 933.28 47.88 ;
   RECT 23.18 47.88 933.28 49.59 ;
   RECT 23.18 49.59 933.28 51.3 ;
   RECT 23.18 51.3 933.28 53.01 ;
   RECT 23.18 53.01 933.28 54.72 ;
   RECT 23.18 54.72 933.28 56.43 ;
   RECT 23.18 56.43 933.28 58.14 ;
   RECT 23.18 58.14 933.28 59.85 ;
   RECT 23.18 59.85 933.28 61.56 ;
   RECT 23.18 61.56 933.28 63.27 ;
   RECT 23.18 63.27 933.28 64.98 ;
   RECT 23.18 64.98 933.28 66.69 ;
   RECT 23.18 66.69 933.28 68.4 ;
   RECT 23.18 68.4 933.28 70.11 ;
   RECT 23.18 70.11 933.28 71.82 ;
   RECT 23.18 71.82 933.28 73.53 ;
   RECT 23.18 73.53 933.28 75.24 ;
   RECT 23.18 75.24 933.28 76.95 ;
   RECT 23.18 76.95 933.28 78.66 ;
   RECT 23.18 78.66 933.28 80.37 ;
   RECT 23.18 80.37 933.28 82.08 ;
   RECT 23.18 82.08 933.28 83.79 ;
   RECT 23.18 83.79 933.28 85.5 ;
   RECT 23.18 85.5 933.28 87.21 ;
   RECT 23.18 87.21 933.28 88.92 ;
   RECT 23.18 88.92 933.28 90.63 ;
   RECT 23.18 90.63 933.28 92.34 ;
   RECT 23.18 92.34 933.28 94.05 ;
   RECT 23.18 94.05 933.28 95.76 ;
   RECT 23.18 95.76 933.28 97.47 ;
   RECT 23.18 97.47 933.28 99.18 ;
   RECT 23.18 99.18 933.28 100.89 ;
   RECT 23.18 100.89 933.28 102.6 ;
   RECT 23.18 102.6 933.28 104.31 ;
   RECT 23.18 104.31 933.28 106.02 ;
   RECT 23.18 106.02 933.28 107.73 ;
   RECT 23.18 107.73 933.28 109.44 ;
   RECT 23.18 109.44 933.28 111.15 ;
   RECT 23.18 111.15 933.28 112.86 ;
   RECT 23.18 112.86 933.28 114.57 ;
   RECT 23.18 114.57 933.28 116.28 ;
   RECT 23.18 116.28 933.28 117.99 ;
   RECT 23.18 117.99 933.28 119.7 ;
   RECT 23.18 119.7 933.28 121.41 ;
   RECT 23.18 121.41 933.28 123.12 ;
   RECT 23.18 123.12 933.28 124.83 ;
   RECT 23.18 124.83 933.28 126.54 ;
   RECT 23.18 126.54 933.28 128.25 ;
   RECT 23.18 128.25 933.28 129.96 ;
   RECT 23.18 129.96 933.28 131.67 ;
   RECT 23.18 131.67 933.28 133.38 ;
   RECT 23.18 133.38 933.28 135.09 ;
   RECT 23.18 135.09 933.28 136.8 ;
   RECT 23.18 136.8 933.28 138.51 ;
   RECT 23.18 138.51 933.28 140.22 ;
   RECT 23.18 140.22 933.28 141.93 ;
   RECT 23.18 141.93 933.28 143.64 ;
   RECT 23.18 143.64 933.28 145.35 ;
   RECT 23.18 145.35 933.28 147.06 ;
   RECT 23.18 147.06 933.28 148.77 ;
   RECT 23.18 148.77 933.28 150.48 ;
   RECT 23.18 150.48 933.28 152.19 ;
   RECT 23.18 152.19 933.28 153.9 ;
   RECT 23.18 153.9 933.28 155.61 ;
   RECT 23.18 155.61 933.28 157.32 ;
   RECT 23.18 157.32 933.28 159.03 ;
   RECT 23.18 159.03 933.28 160.74 ;
   RECT 23.18 160.74 933.28 162.45 ;
   RECT 23.18 162.45 933.28 164.16 ;
   RECT 23.18 164.16 933.28 165.87 ;
   RECT 23.18 165.87 933.28 167.58 ;
   RECT 23.18 167.58 933.28 169.29 ;
   RECT 23.18 169.29 933.28 171.0 ;
   RECT 23.18 171.0 933.28 172.71 ;
   RECT 23.18 172.71 933.28 174.42 ;
   RECT 23.18 174.42 933.28 176.13 ;
   RECT 23.18 176.13 933.28 177.84 ;
   RECT 23.18 177.84 933.28 179.55 ;
   RECT 23.18 179.55 933.28 181.26 ;
   RECT 23.18 181.26 933.28 182.97 ;
   RECT 23.18 182.97 933.28 184.68 ;
   RECT 23.18 184.68 933.28 186.39 ;
   RECT 23.18 186.39 933.28 188.1 ;
   RECT 23.18 188.1 933.28 189.81 ;
   RECT 23.18 189.81 933.28 191.52 ;
   RECT 23.18 191.52 933.28 193.23 ;
   RECT 23.18 193.23 933.28 194.94 ;
   RECT 23.18 194.94 933.28 196.65 ;
   RECT 23.18 196.65 933.28 198.36 ;
   RECT 23.18 198.36 933.28 200.07 ;
   RECT 23.18 200.07 933.28 201.78 ;
   RECT 23.18 201.78 933.28 203.49 ;
   RECT 23.18 203.49 933.28 205.2 ;
   RECT 23.18 205.2 933.28 206.91 ;
   RECT 23.18 206.91 933.28 208.62 ;
   RECT 23.18 208.62 933.28 210.33 ;
   RECT 23.18 210.33 933.28 212.04 ;
   RECT 23.18 212.04 933.28 213.75 ;
   RECT 23.18 213.75 933.28 215.46 ;
   RECT 23.18 215.46 933.28 217.17 ;
   RECT 23.18 217.17 933.28 218.88 ;
   RECT 23.18 218.88 933.28 220.59 ;
   RECT 23.18 220.59 933.28 222.3 ;
   RECT 23.18 222.3 933.28 224.01 ;
   RECT 23.18 224.01 933.28 225.72 ;
   RECT 23.18 225.72 933.28 227.43 ;
   RECT 23.18 227.43 933.28 229.14 ;
   RECT 23.18 229.14 933.28 230.85 ;
   RECT 23.18 230.85 933.28 232.56 ;
   RECT 23.18 232.56 933.28 234.27 ;
   RECT 23.18 234.27 933.28 235.98 ;
   RECT 23.18 235.98 933.28 237.69 ;
   RECT 23.18 237.69 933.28 239.4 ;
   RECT 23.18 239.4 933.28 241.11 ;
   RECT 23.18 241.11 933.28 242.82 ;
   RECT 23.18 242.82 933.28 244.53 ;
   RECT 23.18 244.53 933.28 246.24 ;
   RECT 23.18 246.24 933.28 247.95 ;
   RECT 23.18 247.95 933.28 249.66 ;
   RECT 23.18 249.66 933.28 251.37 ;
   RECT 23.18 251.37 933.28 253.08 ;
   RECT 23.18 253.08 933.28 254.79 ;
   RECT 23.18 254.79 933.28 256.5 ;
   RECT 23.18 256.5 933.28 258.21 ;
   RECT 23.18 258.21 933.28 259.92 ;
   RECT 23.18 259.92 933.28 261.63 ;
   RECT 23.18 261.63 933.28 263.34 ;
   RECT 23.18 263.34 933.28 265.05 ;
   RECT 23.18 265.05 933.28 266.76 ;
   RECT 23.18 266.76 933.28 268.47 ;
   RECT 23.18 268.47 933.28 270.18 ;
   RECT 23.18 270.18 933.28 271.89 ;
   RECT 23.18 271.89 933.28 273.6 ;
   RECT 23.18 273.6 933.28 275.31 ;
   RECT 23.18 275.31 933.28 277.02 ;
   RECT 23.18 277.02 933.28 278.73 ;
   RECT 23.18 278.73 933.28 280.44 ;
   RECT 23.18 280.44 933.28 282.15 ;
   RECT 23.18 282.15 933.28 283.86 ;
   RECT 23.18 283.86 933.28 285.57 ;
   RECT 23.18 285.57 933.28 287.28 ;
   RECT 23.18 287.28 933.28 288.99 ;
   RECT 23.18 288.99 933.28 290.7 ;
   RECT 23.18 290.7 933.28 292.41 ;
   RECT 23.18 292.41 933.28 294.12 ;
   RECT 23.18 294.12 933.28 295.83 ;
   RECT 23.18 295.83 933.28 297.54 ;
   RECT 23.18 297.54 933.28 299.25 ;
   RECT 23.18 299.25 933.28 300.96 ;
   RECT 23.18 300.96 933.28 302.67 ;
   RECT 23.18 302.67 933.28 304.38 ;
   RECT 23.18 304.38 933.28 306.09 ;
   RECT 23.18 306.09 933.28 307.8 ;
   RECT 23.18 307.8 933.28 309.51 ;
   RECT 23.18 309.51 933.28 311.22 ;
   RECT 23.18 311.22 933.28 312.93 ;
   RECT 23.18 312.93 933.28 314.64 ;
   RECT 23.18 314.64 933.28 316.35 ;
   RECT 23.18 316.35 933.28 318.06 ;
   RECT 23.18 318.06 933.28 319.77 ;
   RECT 23.18 319.77 933.28 321.48 ;
   RECT 23.18 321.48 933.28 323.19 ;
   RECT 23.18 323.19 933.28 324.9 ;
   RECT 23.18 324.9 933.28 326.61 ;
   RECT 23.18 326.61 933.28 328.32 ;
   RECT 23.18 328.32 933.28 330.03 ;
   RECT 23.18 330.03 933.28 331.74 ;
   RECT 23.18 331.74 933.28 333.45 ;
   RECT 23.18 333.45 933.28 335.16 ;
   RECT 23.18 335.16 933.28 336.87 ;
   RECT 23.18 336.87 933.28 338.58 ;
   RECT 23.18 338.58 933.28 340.29 ;
   RECT 23.18 340.29 933.28 342.0 ;
   RECT 23.18 342.0 933.28 343.71 ;
   RECT 23.18 343.71 933.28 345.42 ;
   RECT 23.18 345.42 933.28 347.13 ;
   RECT 23.18 347.13 933.28 348.84 ;
   RECT 23.18 348.84 933.28 350.55 ;
   RECT 23.18 350.55 933.28 352.26 ;
   RECT 23.18 352.26 933.28 353.97 ;
   RECT 23.18 353.97 933.28 355.68 ;
   RECT 23.18 355.68 933.28 357.39 ;
   RECT 23.18 357.39 933.28 359.1 ;
   RECT 23.18 359.1 933.28 360.81 ;
   RECT 23.18 360.81 933.28 362.52 ;
   RECT 23.18 362.52 933.28 364.23 ;
   RECT 23.18 364.23 933.28 365.94 ;
   RECT 23.18 365.94 933.28 367.65 ;
   RECT 23.18 367.65 933.28 369.36 ;
   RECT 23.18 369.36 933.28 371.07 ;
   RECT 23.18 371.07 933.28 372.78 ;
   RECT 23.18 372.78 933.28 374.49 ;
   RECT 23.18 374.49 933.28 376.2 ;
   RECT 23.18 376.2 933.28 377.91 ;
   RECT 23.18 377.91 933.28 379.62 ;
   RECT 23.18 379.62 933.28 381.33 ;
   RECT 23.18 381.33 933.28 383.04 ;
   RECT 23.18 383.04 933.28 384.75 ;
   RECT 23.18 384.75 933.28 386.46 ;
   RECT 23.18 386.46 933.28 388.17 ;
   RECT 23.18 388.17 933.28 389.88 ;
   RECT 23.18 389.88 933.28 391.59 ;
   RECT 23.18 391.59 933.28 393.3 ;
   RECT 23.18 393.3 933.28 395.01 ;
   RECT 23.18 395.01 933.28 396.72 ;
   RECT 23.18 396.72 933.28 398.43 ;
   RECT 23.18 398.43 933.28 400.14 ;
   RECT 23.18 400.14 933.28 401.85 ;
   RECT 23.18 401.85 933.28 403.56 ;
   RECT 23.18 403.56 933.28 405.27 ;
   RECT 23.18 405.27 933.28 406.98 ;
   RECT 23.18 406.98 933.28 408.69 ;
   RECT 23.18 408.69 933.28 410.4 ;
   RECT 23.18 410.4 933.28 412.11 ;
   RECT 23.18 412.11 933.28 413.82 ;
   RECT 23.18 413.82 933.28 415.53 ;
   RECT 23.18 415.53 933.28 417.24 ;
   RECT 23.18 417.24 933.28 418.95 ;
   RECT 23.18 418.95 933.28 420.66 ;
   RECT 23.18 420.66 933.28 422.37 ;
   RECT 23.18 422.37 933.28 424.08 ;
   RECT 23.18 424.08 933.28 425.79 ;
   RECT 23.18 425.79 933.28 427.5 ;
   RECT 23.18 427.5 933.28 429.21 ;
   RECT 23.18 429.21 933.28 430.92 ;
   RECT 0.0 430.92 933.28 432.63 ;
   RECT 0.0 432.63 933.28 434.34 ;
   RECT 0.0 434.34 933.28 436.05 ;
   RECT 0.0 436.05 933.28 437.76 ;
   RECT 0.0 437.76 933.28 439.47 ;
   RECT 0.0 439.47 933.28 441.18 ;
   RECT 0.0 441.18 933.28 442.89 ;
   RECT 0.0 442.89 933.28 444.6 ;
   RECT 0.0 444.6 933.28 446.31 ;
   RECT 0.0 446.31 933.28 448.02 ;
   RECT 0.0 448.02 933.28 449.73 ;
   RECT 0.0 449.73 933.28 451.44 ;
   RECT 0.0 451.44 933.28 453.15 ;
   RECT 0.0 453.15 933.28 454.86 ;
   RECT 0.0 454.86 933.28 456.57 ;
   RECT 0.0 456.57 933.28 458.28 ;
   RECT 0.0 458.28 933.28 459.99 ;
   RECT 23.18 459.99 933.28 461.7 ;
   RECT 23.18 461.7 933.28 463.41 ;
   RECT 23.18 463.41 933.28 465.12 ;
   RECT 23.18 465.12 933.28 466.83 ;
   RECT 23.18 466.83 933.28 468.54 ;
   RECT 23.18 468.54 933.28 470.25 ;
   RECT 23.18 470.25 933.28 471.96 ;
   RECT 23.18 471.96 933.28 473.67 ;
   RECT 23.18 473.67 933.28 475.38 ;
   RECT 23.18 475.38 933.28 477.09 ;
   RECT 23.18 477.09 933.28 478.8 ;
   RECT 23.18 478.8 933.28 480.51 ;
   RECT 23.18 480.51 933.28 482.22 ;
   RECT 23.18 482.22 933.28 483.93 ;
   RECT 23.18 483.93 933.28 485.64 ;
   RECT 23.18 485.64 933.28 487.35 ;
   RECT 23.18 487.35 933.28 489.06 ;
   RECT 23.18 489.06 933.28 490.77 ;
   RECT 23.18 490.77 933.28 492.48 ;
   RECT 23.18 492.48 933.28 494.19 ;
   RECT 23.18 494.19 933.28 495.9 ;
   RECT 23.18 495.9 933.28 497.61 ;
   RECT 23.18 497.61 933.28 499.32 ;
   RECT 23.18 499.32 933.28 501.03 ;
   RECT 23.18 501.03 933.28 502.74 ;
   RECT 23.18 502.74 933.28 504.45 ;
   RECT 23.18 504.45 933.28 506.16 ;
   RECT 23.18 506.16 933.28 507.87 ;
   RECT 23.18 507.87 933.28 509.58 ;
   RECT 23.18 509.58 933.28 511.29 ;
   RECT 23.18 511.29 933.28 513.0 ;
   RECT 23.18 513.0 933.28 514.71 ;
   RECT 23.18 514.71 933.28 516.42 ;
   RECT 23.18 516.42 933.28 518.13 ;
   RECT 23.18 518.13 933.28 519.84 ;
   RECT 23.18 519.84 933.28 521.55 ;
   RECT 23.18 521.55 933.28 523.26 ;
   RECT 23.18 523.26 933.28 524.97 ;
   RECT 23.18 524.97 933.28 526.68 ;
   RECT 23.18 526.68 933.28 528.39 ;
   RECT 23.18 528.39 933.28 530.1 ;
   RECT 23.18 530.1 933.28 531.81 ;
   RECT 23.18 531.81 933.28 533.52 ;
   RECT 23.18 533.52 933.28 535.23 ;
   RECT 23.18 535.23 933.28 536.94 ;
   RECT 23.18 536.94 933.28 538.65 ;
   RECT 23.18 538.65 933.28 540.36 ;
   RECT 23.18 540.36 933.28 542.07 ;
   RECT 23.18 542.07 933.28 543.78 ;
   RECT 23.18 543.78 933.28 545.49 ;
   RECT 23.18 545.49 933.28 547.2 ;
   RECT 23.18 547.2 933.28 548.91 ;
   RECT 23.18 548.91 933.28 550.62 ;
   RECT 23.18 550.62 933.28 552.33 ;
   RECT 23.18 552.33 933.28 554.04 ;
   RECT 23.18 554.04 933.28 555.75 ;
   RECT 23.18 555.75 933.28 557.46 ;
   RECT 23.18 557.46 933.28 559.17 ;
   RECT 23.18 559.17 933.28 560.88 ;
   RECT 23.18 560.88 933.28 562.59 ;
   RECT 23.18 562.59 933.28 564.3 ;
   RECT 23.18 564.3 933.28 566.01 ;
   RECT 23.18 566.01 933.28 567.72 ;
   RECT 23.18 567.72 933.28 569.43 ;
   RECT 23.18 569.43 933.28 571.14 ;
   RECT 23.18 571.14 933.28 572.85 ;
   RECT 23.18 572.85 933.28 574.56 ;
   RECT 23.18 574.56 933.28 576.27 ;
   RECT 23.18 576.27 933.28 577.98 ;
   RECT 23.18 577.98 933.28 579.69 ;
   RECT 23.18 579.69 933.28 581.4 ;
   RECT 23.18 581.4 933.28 583.11 ;
   RECT 23.18 583.11 933.28 584.82 ;
   RECT 23.18 584.82 933.28 586.53 ;
   RECT 23.18 586.53 933.28 588.24 ;
   RECT 23.18 588.24 933.28 589.95 ;
   RECT 23.18 589.95 933.28 591.66 ;
   RECT 23.18 591.66 933.28 593.37 ;
   RECT 23.18 593.37 933.28 595.08 ;
   RECT 23.18 595.08 933.28 596.79 ;
   RECT 23.18 596.79 933.28 598.5 ;
   RECT 23.18 598.5 933.28 600.21 ;
   RECT 23.18 600.21 933.28 601.92 ;
   RECT 23.18 601.92 933.28 603.63 ;
   RECT 23.18 603.63 933.28 605.34 ;
   RECT 23.18 605.34 933.28 607.05 ;
   RECT 23.18 607.05 933.28 608.76 ;
   RECT 23.18 608.76 933.28 610.47 ;
   RECT 23.18 610.47 933.28 612.18 ;
   RECT 23.18 612.18 933.28 613.89 ;
   RECT 23.18 613.89 933.28 615.6 ;
   RECT 23.18 615.6 933.28 617.31 ;
   RECT 23.18 617.31 933.28 619.02 ;
   RECT 23.18 619.02 933.28 620.73 ;
   RECT 23.18 620.73 933.28 622.44 ;
   RECT 23.18 622.44 933.28 624.15 ;
   RECT 23.18 624.15 933.28 625.86 ;
   RECT 23.18 625.86 933.28 627.57 ;
   RECT 23.18 627.57 933.28 629.28 ;
   RECT 23.18 629.28 933.28 630.99 ;
   RECT 23.18 630.99 933.28 632.7 ;
   RECT 23.18 632.7 933.28 634.41 ;
   RECT 23.18 634.41 933.28 636.12 ;
   RECT 23.18 636.12 933.28 637.83 ;
   RECT 23.18 637.83 933.28 639.54 ;
   RECT 23.18 639.54 933.28 641.25 ;
   RECT 23.18 641.25 933.28 642.96 ;
   RECT 23.18 642.96 933.28 644.67 ;
   RECT 23.18 644.67 933.28 646.38 ;
   RECT 23.18 646.38 933.28 648.09 ;
   RECT 23.18 648.09 933.28 649.8 ;
   RECT 23.18 649.8 933.28 651.51 ;
   RECT 23.18 651.51 933.28 653.22 ;
   RECT 23.18 653.22 933.28 654.93 ;
   RECT 23.18 654.93 933.28 656.64 ;
   RECT 23.18 656.64 933.28 658.35 ;
   RECT 23.18 658.35 933.28 660.06 ;
   RECT 23.18 660.06 933.28 661.77 ;
   RECT 23.18 661.77 933.28 663.48 ;
   RECT 23.18 663.48 933.28 665.19 ;
   RECT 23.18 665.19 933.28 666.9 ;
   RECT 23.18 666.9 933.28 668.61 ;
   RECT 23.18 668.61 933.28 670.32 ;
   RECT 23.18 670.32 933.28 672.03 ;
   RECT 23.18 672.03 933.28 673.74 ;
   RECT 23.18 673.74 933.28 675.45 ;
   RECT 23.18 675.45 933.28 677.16 ;
   RECT 23.18 677.16 933.28 678.87 ;
   RECT 23.18 678.87 933.28 680.58 ;
   RECT 23.18 680.58 933.28 682.29 ;
   RECT 23.18 682.29 933.28 684.0 ;
   RECT 23.18 684.0 933.28 685.71 ;
   RECT 23.18 685.71 933.28 687.42 ;
   RECT 23.18 687.42 933.28 689.13 ;
   RECT 23.18 689.13 933.28 690.84 ;
   RECT 23.18 690.84 933.28 692.55 ;
   RECT 23.18 692.55 933.28 694.26 ;
   RECT 23.18 694.26 933.28 695.97 ;
   RECT 23.18 695.97 933.28 697.68 ;
   RECT 23.18 697.68 933.28 699.39 ;
   RECT 23.18 699.39 933.28 701.1 ;
   RECT 23.18 701.1 933.28 702.81 ;
   RECT 23.18 702.81 933.28 704.52 ;
   RECT 23.18 704.52 933.28 706.23 ;
   RECT 23.18 706.23 933.28 707.94 ;
   RECT 23.18 707.94 933.28 709.65 ;
   RECT 23.18 709.65 933.28 711.36 ;
   RECT 23.18 711.36 933.28 713.07 ;
   RECT 23.18 713.07 933.28 714.78 ;
   RECT 23.18 714.78 933.28 716.49 ;
   RECT 23.18 716.49 933.28 718.2 ;
   RECT 23.18 718.2 933.28 719.91 ;
   RECT 23.18 719.91 933.28 721.62 ;
   RECT 23.18 721.62 933.28 723.33 ;
   RECT 23.18 723.33 933.28 725.04 ;
   RECT 23.18 725.04 933.28 726.75 ;
   RECT 23.18 726.75 933.28 728.46 ;
   RECT 23.18 728.46 933.28 730.17 ;
   RECT 23.18 730.17 933.28 731.88 ;
   RECT 23.18 731.88 933.28 733.59 ;
   RECT 23.18 733.59 933.28 735.3 ;
   RECT 23.18 735.3 933.28 737.01 ;
   RECT 23.18 737.01 933.28 738.72 ;
   RECT 23.18 738.72 933.28 740.43 ;
   RECT 23.18 740.43 933.28 742.14 ;
   RECT 23.18 742.14 933.28 743.85 ;
   RECT 23.18 743.85 933.28 745.56 ;
   RECT 23.18 745.56 933.28 747.27 ;
   RECT 23.18 747.27 933.28 748.98 ;
   RECT 23.18 748.98 933.28 750.69 ;
   RECT 23.18 750.69 933.28 752.4 ;
   RECT 23.18 752.4 933.28 754.11 ;
   RECT 23.18 754.11 933.28 755.82 ;
   RECT 23.18 755.82 933.28 757.53 ;
   RECT 23.18 757.53 933.28 759.24 ;
   RECT 23.18 759.24 933.28 760.95 ;
   RECT 23.18 760.95 933.28 762.66 ;
   RECT 23.18 762.66 933.28 764.37 ;
   RECT 23.18 764.37 933.28 766.08 ;
   RECT 23.18 766.08 933.28 767.79 ;
   RECT 23.18 767.79 933.28 769.5 ;
   RECT 23.18 769.5 933.28 771.21 ;
   RECT 23.18 771.21 933.28 772.92 ;
   RECT 23.18 772.92 933.28 774.63 ;
   RECT 23.18 774.63 933.28 776.34 ;
   RECT 23.18 776.34 933.28 778.05 ;
   RECT 23.18 778.05 933.28 779.76 ;
   RECT 23.18 779.76 933.28 781.47 ;
   RECT 23.18 781.47 933.28 783.18 ;
   RECT 23.18 783.18 933.28 784.89 ;
   RECT 23.18 784.89 933.28 786.6 ;
   RECT 23.18 786.6 933.28 788.31 ;
   RECT 23.18 788.31 933.28 790.02 ;
   RECT 23.18 790.02 933.28 791.73 ;
   RECT 23.18 791.73 933.28 793.44 ;
   RECT 23.18 793.44 933.28 795.15 ;
   RECT 23.18 795.15 933.28 796.86 ;
   RECT 23.18 796.86 933.28 798.57 ;
   RECT 23.18 798.57 933.28 800.28 ;
   RECT 23.18 800.28 933.28 801.99 ;
   RECT 23.18 801.99 933.28 803.7 ;
   RECT 23.18 803.7 933.28 805.41 ;
   RECT 23.18 805.41 933.28 807.12 ;
   RECT 23.18 807.12 933.28 808.83 ;
   RECT 23.18 808.83 933.28 810.54 ;
   RECT 23.18 810.54 933.28 812.25 ;
   RECT 23.18 812.25 933.28 813.96 ;
   RECT 23.18 813.96 933.28 815.67 ;
   RECT 23.18 815.67 933.28 817.38 ;
   RECT 23.18 817.38 933.28 819.09 ;
   RECT 23.18 819.09 933.28 820.8 ;
   RECT 23.18 820.8 933.28 822.51 ;
   RECT 23.18 822.51 933.28 824.22 ;
   RECT 23.18 824.22 933.28 825.93 ;
   RECT 23.18 825.93 933.28 827.64 ;
   RECT 23.18 827.64 933.28 829.35 ;
   RECT 23.18 829.35 933.28 831.06 ;
   RECT 23.18 831.06 933.28 832.77 ;
   RECT 23.18 832.77 933.28 834.48 ;
   RECT 23.18 834.48 933.28 836.19 ;
   RECT 23.18 836.19 933.28 837.9 ;
   RECT 23.18 837.9 933.28 839.61 ;
   RECT 23.18 839.61 933.28 841.32 ;
   RECT 23.18 841.32 933.28 843.03 ;
   RECT 23.18 843.03 933.28 844.74 ;
   RECT 23.18 844.74 933.28 846.45 ;
   RECT 23.18 846.45 933.28 848.16 ;
   RECT 23.18 848.16 933.28 849.87 ;
   RECT 23.18 849.87 933.28 851.58 ;
   RECT 23.18 851.58 933.28 853.29 ;
   RECT 23.18 853.29 933.28 855.0 ;
   RECT 23.18 855.0 933.28 856.71 ;
   RECT 23.18 856.71 933.28 858.42 ;
   RECT 23.18 858.42 933.28 860.13 ;
   RECT 23.18 860.13 933.28 861.84 ;
   RECT 23.18 861.84 933.28 863.55 ;
   RECT 23.18 863.55 933.28 865.26 ;
   RECT 23.18 865.26 933.28 866.97 ;
   RECT 23.18 866.97 933.28 868.68 ;
   RECT 23.18 868.68 933.28 870.39 ;
   RECT 23.18 870.39 933.28 872.1 ;
   RECT 23.18 872.1 933.28 873.81 ;
   RECT 23.18 873.81 933.28 875.52 ;
   RECT 23.18 875.52 933.28 877.23 ;
   RECT 23.18 877.23 933.28 878.94 ;
  LAYER via3 ;
   RECT 23.18 0.0 933.28 1.71 ;
   RECT 23.18 1.71 933.28 3.42 ;
   RECT 23.18 3.42 933.28 5.13 ;
   RECT 23.18 5.13 933.28 6.84 ;
   RECT 23.18 6.84 933.28 8.55 ;
   RECT 23.18 8.55 933.28 10.26 ;
   RECT 23.18 10.26 933.28 11.97 ;
   RECT 23.18 11.97 933.28 13.68 ;
   RECT 23.18 13.68 933.28 15.39 ;
   RECT 23.18 15.39 933.28 17.1 ;
   RECT 23.18 17.1 933.28 18.81 ;
   RECT 23.18 18.81 933.28 20.52 ;
   RECT 23.18 20.52 933.28 22.23 ;
   RECT 23.18 22.23 933.28 23.94 ;
   RECT 23.18 23.94 933.28 25.65 ;
   RECT 23.18 25.65 933.28 27.36 ;
   RECT 23.18 27.36 933.28 29.07 ;
   RECT 23.18 29.07 933.28 30.78 ;
   RECT 23.18 30.78 933.28 32.49 ;
   RECT 23.18 32.49 933.28 34.2 ;
   RECT 23.18 34.2 933.28 35.91 ;
   RECT 23.18 35.91 933.28 37.62 ;
   RECT 23.18 37.62 933.28 39.33 ;
   RECT 23.18 39.33 933.28 41.04 ;
   RECT 23.18 41.04 933.28 42.75 ;
   RECT 23.18 42.75 933.28 44.46 ;
   RECT 23.18 44.46 933.28 46.17 ;
   RECT 23.18 46.17 933.28 47.88 ;
   RECT 23.18 47.88 933.28 49.59 ;
   RECT 23.18 49.59 933.28 51.3 ;
   RECT 23.18 51.3 933.28 53.01 ;
   RECT 23.18 53.01 933.28 54.72 ;
   RECT 23.18 54.72 933.28 56.43 ;
   RECT 23.18 56.43 933.28 58.14 ;
   RECT 23.18 58.14 933.28 59.85 ;
   RECT 23.18 59.85 933.28 61.56 ;
   RECT 23.18 61.56 933.28 63.27 ;
   RECT 23.18 63.27 933.28 64.98 ;
   RECT 23.18 64.98 933.28 66.69 ;
   RECT 23.18 66.69 933.28 68.4 ;
   RECT 23.18 68.4 933.28 70.11 ;
   RECT 23.18 70.11 933.28 71.82 ;
   RECT 23.18 71.82 933.28 73.53 ;
   RECT 23.18 73.53 933.28 75.24 ;
   RECT 23.18 75.24 933.28 76.95 ;
   RECT 23.18 76.95 933.28 78.66 ;
   RECT 23.18 78.66 933.28 80.37 ;
   RECT 23.18 80.37 933.28 82.08 ;
   RECT 23.18 82.08 933.28 83.79 ;
   RECT 23.18 83.79 933.28 85.5 ;
   RECT 23.18 85.5 933.28 87.21 ;
   RECT 23.18 87.21 933.28 88.92 ;
   RECT 23.18 88.92 933.28 90.63 ;
   RECT 23.18 90.63 933.28 92.34 ;
   RECT 23.18 92.34 933.28 94.05 ;
   RECT 23.18 94.05 933.28 95.76 ;
   RECT 23.18 95.76 933.28 97.47 ;
   RECT 23.18 97.47 933.28 99.18 ;
   RECT 23.18 99.18 933.28 100.89 ;
   RECT 23.18 100.89 933.28 102.6 ;
   RECT 23.18 102.6 933.28 104.31 ;
   RECT 23.18 104.31 933.28 106.02 ;
   RECT 23.18 106.02 933.28 107.73 ;
   RECT 23.18 107.73 933.28 109.44 ;
   RECT 23.18 109.44 933.28 111.15 ;
   RECT 23.18 111.15 933.28 112.86 ;
   RECT 23.18 112.86 933.28 114.57 ;
   RECT 23.18 114.57 933.28 116.28 ;
   RECT 23.18 116.28 933.28 117.99 ;
   RECT 23.18 117.99 933.28 119.7 ;
   RECT 23.18 119.7 933.28 121.41 ;
   RECT 23.18 121.41 933.28 123.12 ;
   RECT 23.18 123.12 933.28 124.83 ;
   RECT 23.18 124.83 933.28 126.54 ;
   RECT 23.18 126.54 933.28 128.25 ;
   RECT 23.18 128.25 933.28 129.96 ;
   RECT 23.18 129.96 933.28 131.67 ;
   RECT 23.18 131.67 933.28 133.38 ;
   RECT 23.18 133.38 933.28 135.09 ;
   RECT 23.18 135.09 933.28 136.8 ;
   RECT 23.18 136.8 933.28 138.51 ;
   RECT 23.18 138.51 933.28 140.22 ;
   RECT 23.18 140.22 933.28 141.93 ;
   RECT 23.18 141.93 933.28 143.64 ;
   RECT 23.18 143.64 933.28 145.35 ;
   RECT 23.18 145.35 933.28 147.06 ;
   RECT 23.18 147.06 933.28 148.77 ;
   RECT 23.18 148.77 933.28 150.48 ;
   RECT 23.18 150.48 933.28 152.19 ;
   RECT 23.18 152.19 933.28 153.9 ;
   RECT 23.18 153.9 933.28 155.61 ;
   RECT 23.18 155.61 933.28 157.32 ;
   RECT 23.18 157.32 933.28 159.03 ;
   RECT 23.18 159.03 933.28 160.74 ;
   RECT 23.18 160.74 933.28 162.45 ;
   RECT 23.18 162.45 933.28 164.16 ;
   RECT 23.18 164.16 933.28 165.87 ;
   RECT 23.18 165.87 933.28 167.58 ;
   RECT 23.18 167.58 933.28 169.29 ;
   RECT 23.18 169.29 933.28 171.0 ;
   RECT 23.18 171.0 933.28 172.71 ;
   RECT 23.18 172.71 933.28 174.42 ;
   RECT 23.18 174.42 933.28 176.13 ;
   RECT 23.18 176.13 933.28 177.84 ;
   RECT 23.18 177.84 933.28 179.55 ;
   RECT 23.18 179.55 933.28 181.26 ;
   RECT 23.18 181.26 933.28 182.97 ;
   RECT 23.18 182.97 933.28 184.68 ;
   RECT 23.18 184.68 933.28 186.39 ;
   RECT 23.18 186.39 933.28 188.1 ;
   RECT 23.18 188.1 933.28 189.81 ;
   RECT 23.18 189.81 933.28 191.52 ;
   RECT 23.18 191.52 933.28 193.23 ;
   RECT 23.18 193.23 933.28 194.94 ;
   RECT 23.18 194.94 933.28 196.65 ;
   RECT 23.18 196.65 933.28 198.36 ;
   RECT 23.18 198.36 933.28 200.07 ;
   RECT 23.18 200.07 933.28 201.78 ;
   RECT 23.18 201.78 933.28 203.49 ;
   RECT 23.18 203.49 933.28 205.2 ;
   RECT 23.18 205.2 933.28 206.91 ;
   RECT 23.18 206.91 933.28 208.62 ;
   RECT 23.18 208.62 933.28 210.33 ;
   RECT 23.18 210.33 933.28 212.04 ;
   RECT 23.18 212.04 933.28 213.75 ;
   RECT 23.18 213.75 933.28 215.46 ;
   RECT 23.18 215.46 933.28 217.17 ;
   RECT 23.18 217.17 933.28 218.88 ;
   RECT 23.18 218.88 933.28 220.59 ;
   RECT 23.18 220.59 933.28 222.3 ;
   RECT 23.18 222.3 933.28 224.01 ;
   RECT 23.18 224.01 933.28 225.72 ;
   RECT 23.18 225.72 933.28 227.43 ;
   RECT 23.18 227.43 933.28 229.14 ;
   RECT 23.18 229.14 933.28 230.85 ;
   RECT 23.18 230.85 933.28 232.56 ;
   RECT 23.18 232.56 933.28 234.27 ;
   RECT 23.18 234.27 933.28 235.98 ;
   RECT 23.18 235.98 933.28 237.69 ;
   RECT 23.18 237.69 933.28 239.4 ;
   RECT 23.18 239.4 933.28 241.11 ;
   RECT 23.18 241.11 933.28 242.82 ;
   RECT 23.18 242.82 933.28 244.53 ;
   RECT 23.18 244.53 933.28 246.24 ;
   RECT 23.18 246.24 933.28 247.95 ;
   RECT 23.18 247.95 933.28 249.66 ;
   RECT 23.18 249.66 933.28 251.37 ;
   RECT 23.18 251.37 933.28 253.08 ;
   RECT 23.18 253.08 933.28 254.79 ;
   RECT 23.18 254.79 933.28 256.5 ;
   RECT 23.18 256.5 933.28 258.21 ;
   RECT 23.18 258.21 933.28 259.92 ;
   RECT 23.18 259.92 933.28 261.63 ;
   RECT 23.18 261.63 933.28 263.34 ;
   RECT 23.18 263.34 933.28 265.05 ;
   RECT 23.18 265.05 933.28 266.76 ;
   RECT 23.18 266.76 933.28 268.47 ;
   RECT 23.18 268.47 933.28 270.18 ;
   RECT 23.18 270.18 933.28 271.89 ;
   RECT 23.18 271.89 933.28 273.6 ;
   RECT 23.18 273.6 933.28 275.31 ;
   RECT 23.18 275.31 933.28 277.02 ;
   RECT 23.18 277.02 933.28 278.73 ;
   RECT 23.18 278.73 933.28 280.44 ;
   RECT 23.18 280.44 933.28 282.15 ;
   RECT 23.18 282.15 933.28 283.86 ;
   RECT 23.18 283.86 933.28 285.57 ;
   RECT 23.18 285.57 933.28 287.28 ;
   RECT 23.18 287.28 933.28 288.99 ;
   RECT 23.18 288.99 933.28 290.7 ;
   RECT 23.18 290.7 933.28 292.41 ;
   RECT 23.18 292.41 933.28 294.12 ;
   RECT 23.18 294.12 933.28 295.83 ;
   RECT 23.18 295.83 933.28 297.54 ;
   RECT 23.18 297.54 933.28 299.25 ;
   RECT 23.18 299.25 933.28 300.96 ;
   RECT 23.18 300.96 933.28 302.67 ;
   RECT 23.18 302.67 933.28 304.38 ;
   RECT 23.18 304.38 933.28 306.09 ;
   RECT 23.18 306.09 933.28 307.8 ;
   RECT 23.18 307.8 933.28 309.51 ;
   RECT 23.18 309.51 933.28 311.22 ;
   RECT 23.18 311.22 933.28 312.93 ;
   RECT 23.18 312.93 933.28 314.64 ;
   RECT 23.18 314.64 933.28 316.35 ;
   RECT 23.18 316.35 933.28 318.06 ;
   RECT 23.18 318.06 933.28 319.77 ;
   RECT 23.18 319.77 933.28 321.48 ;
   RECT 23.18 321.48 933.28 323.19 ;
   RECT 23.18 323.19 933.28 324.9 ;
   RECT 23.18 324.9 933.28 326.61 ;
   RECT 23.18 326.61 933.28 328.32 ;
   RECT 23.18 328.32 933.28 330.03 ;
   RECT 23.18 330.03 933.28 331.74 ;
   RECT 23.18 331.74 933.28 333.45 ;
   RECT 23.18 333.45 933.28 335.16 ;
   RECT 23.18 335.16 933.28 336.87 ;
   RECT 23.18 336.87 933.28 338.58 ;
   RECT 23.18 338.58 933.28 340.29 ;
   RECT 23.18 340.29 933.28 342.0 ;
   RECT 23.18 342.0 933.28 343.71 ;
   RECT 23.18 343.71 933.28 345.42 ;
   RECT 23.18 345.42 933.28 347.13 ;
   RECT 23.18 347.13 933.28 348.84 ;
   RECT 23.18 348.84 933.28 350.55 ;
   RECT 23.18 350.55 933.28 352.26 ;
   RECT 23.18 352.26 933.28 353.97 ;
   RECT 23.18 353.97 933.28 355.68 ;
   RECT 23.18 355.68 933.28 357.39 ;
   RECT 23.18 357.39 933.28 359.1 ;
   RECT 23.18 359.1 933.28 360.81 ;
   RECT 23.18 360.81 933.28 362.52 ;
   RECT 23.18 362.52 933.28 364.23 ;
   RECT 23.18 364.23 933.28 365.94 ;
   RECT 23.18 365.94 933.28 367.65 ;
   RECT 23.18 367.65 933.28 369.36 ;
   RECT 23.18 369.36 933.28 371.07 ;
   RECT 23.18 371.07 933.28 372.78 ;
   RECT 23.18 372.78 933.28 374.49 ;
   RECT 23.18 374.49 933.28 376.2 ;
   RECT 23.18 376.2 933.28 377.91 ;
   RECT 23.18 377.91 933.28 379.62 ;
   RECT 23.18 379.62 933.28 381.33 ;
   RECT 23.18 381.33 933.28 383.04 ;
   RECT 23.18 383.04 933.28 384.75 ;
   RECT 23.18 384.75 933.28 386.46 ;
   RECT 23.18 386.46 933.28 388.17 ;
   RECT 23.18 388.17 933.28 389.88 ;
   RECT 23.18 389.88 933.28 391.59 ;
   RECT 23.18 391.59 933.28 393.3 ;
   RECT 23.18 393.3 933.28 395.01 ;
   RECT 23.18 395.01 933.28 396.72 ;
   RECT 23.18 396.72 933.28 398.43 ;
   RECT 23.18 398.43 933.28 400.14 ;
   RECT 23.18 400.14 933.28 401.85 ;
   RECT 23.18 401.85 933.28 403.56 ;
   RECT 23.18 403.56 933.28 405.27 ;
   RECT 23.18 405.27 933.28 406.98 ;
   RECT 23.18 406.98 933.28 408.69 ;
   RECT 23.18 408.69 933.28 410.4 ;
   RECT 23.18 410.4 933.28 412.11 ;
   RECT 23.18 412.11 933.28 413.82 ;
   RECT 23.18 413.82 933.28 415.53 ;
   RECT 23.18 415.53 933.28 417.24 ;
   RECT 23.18 417.24 933.28 418.95 ;
   RECT 23.18 418.95 933.28 420.66 ;
   RECT 23.18 420.66 933.28 422.37 ;
   RECT 23.18 422.37 933.28 424.08 ;
   RECT 23.18 424.08 933.28 425.79 ;
   RECT 23.18 425.79 933.28 427.5 ;
   RECT 23.18 427.5 933.28 429.21 ;
   RECT 23.18 429.21 933.28 430.92 ;
   RECT 0.0 430.92 933.28 432.63 ;
   RECT 0.0 432.63 933.28 434.34 ;
   RECT 0.0 434.34 933.28 436.05 ;
   RECT 0.0 436.05 933.28 437.76 ;
   RECT 0.0 437.76 933.28 439.47 ;
   RECT 0.0 439.47 933.28 441.18 ;
   RECT 0.0 441.18 933.28 442.89 ;
   RECT 0.0 442.89 933.28 444.6 ;
   RECT 0.0 444.6 933.28 446.31 ;
   RECT 0.0 446.31 933.28 448.02 ;
   RECT 0.0 448.02 933.28 449.73 ;
   RECT 0.0 449.73 933.28 451.44 ;
   RECT 0.0 451.44 933.28 453.15 ;
   RECT 0.0 453.15 933.28 454.86 ;
   RECT 0.0 454.86 933.28 456.57 ;
   RECT 0.0 456.57 933.28 458.28 ;
   RECT 0.0 458.28 933.28 459.99 ;
   RECT 23.18 459.99 933.28 461.7 ;
   RECT 23.18 461.7 933.28 463.41 ;
   RECT 23.18 463.41 933.28 465.12 ;
   RECT 23.18 465.12 933.28 466.83 ;
   RECT 23.18 466.83 933.28 468.54 ;
   RECT 23.18 468.54 933.28 470.25 ;
   RECT 23.18 470.25 933.28 471.96 ;
   RECT 23.18 471.96 933.28 473.67 ;
   RECT 23.18 473.67 933.28 475.38 ;
   RECT 23.18 475.38 933.28 477.09 ;
   RECT 23.18 477.09 933.28 478.8 ;
   RECT 23.18 478.8 933.28 480.51 ;
   RECT 23.18 480.51 933.28 482.22 ;
   RECT 23.18 482.22 933.28 483.93 ;
   RECT 23.18 483.93 933.28 485.64 ;
   RECT 23.18 485.64 933.28 487.35 ;
   RECT 23.18 487.35 933.28 489.06 ;
   RECT 23.18 489.06 933.28 490.77 ;
   RECT 23.18 490.77 933.28 492.48 ;
   RECT 23.18 492.48 933.28 494.19 ;
   RECT 23.18 494.19 933.28 495.9 ;
   RECT 23.18 495.9 933.28 497.61 ;
   RECT 23.18 497.61 933.28 499.32 ;
   RECT 23.18 499.32 933.28 501.03 ;
   RECT 23.18 501.03 933.28 502.74 ;
   RECT 23.18 502.74 933.28 504.45 ;
   RECT 23.18 504.45 933.28 506.16 ;
   RECT 23.18 506.16 933.28 507.87 ;
   RECT 23.18 507.87 933.28 509.58 ;
   RECT 23.18 509.58 933.28 511.29 ;
   RECT 23.18 511.29 933.28 513.0 ;
   RECT 23.18 513.0 933.28 514.71 ;
   RECT 23.18 514.71 933.28 516.42 ;
   RECT 23.18 516.42 933.28 518.13 ;
   RECT 23.18 518.13 933.28 519.84 ;
   RECT 23.18 519.84 933.28 521.55 ;
   RECT 23.18 521.55 933.28 523.26 ;
   RECT 23.18 523.26 933.28 524.97 ;
   RECT 23.18 524.97 933.28 526.68 ;
   RECT 23.18 526.68 933.28 528.39 ;
   RECT 23.18 528.39 933.28 530.1 ;
   RECT 23.18 530.1 933.28 531.81 ;
   RECT 23.18 531.81 933.28 533.52 ;
   RECT 23.18 533.52 933.28 535.23 ;
   RECT 23.18 535.23 933.28 536.94 ;
   RECT 23.18 536.94 933.28 538.65 ;
   RECT 23.18 538.65 933.28 540.36 ;
   RECT 23.18 540.36 933.28 542.07 ;
   RECT 23.18 542.07 933.28 543.78 ;
   RECT 23.18 543.78 933.28 545.49 ;
   RECT 23.18 545.49 933.28 547.2 ;
   RECT 23.18 547.2 933.28 548.91 ;
   RECT 23.18 548.91 933.28 550.62 ;
   RECT 23.18 550.62 933.28 552.33 ;
   RECT 23.18 552.33 933.28 554.04 ;
   RECT 23.18 554.04 933.28 555.75 ;
   RECT 23.18 555.75 933.28 557.46 ;
   RECT 23.18 557.46 933.28 559.17 ;
   RECT 23.18 559.17 933.28 560.88 ;
   RECT 23.18 560.88 933.28 562.59 ;
   RECT 23.18 562.59 933.28 564.3 ;
   RECT 23.18 564.3 933.28 566.01 ;
   RECT 23.18 566.01 933.28 567.72 ;
   RECT 23.18 567.72 933.28 569.43 ;
   RECT 23.18 569.43 933.28 571.14 ;
   RECT 23.18 571.14 933.28 572.85 ;
   RECT 23.18 572.85 933.28 574.56 ;
   RECT 23.18 574.56 933.28 576.27 ;
   RECT 23.18 576.27 933.28 577.98 ;
   RECT 23.18 577.98 933.28 579.69 ;
   RECT 23.18 579.69 933.28 581.4 ;
   RECT 23.18 581.4 933.28 583.11 ;
   RECT 23.18 583.11 933.28 584.82 ;
   RECT 23.18 584.82 933.28 586.53 ;
   RECT 23.18 586.53 933.28 588.24 ;
   RECT 23.18 588.24 933.28 589.95 ;
   RECT 23.18 589.95 933.28 591.66 ;
   RECT 23.18 591.66 933.28 593.37 ;
   RECT 23.18 593.37 933.28 595.08 ;
   RECT 23.18 595.08 933.28 596.79 ;
   RECT 23.18 596.79 933.28 598.5 ;
   RECT 23.18 598.5 933.28 600.21 ;
   RECT 23.18 600.21 933.28 601.92 ;
   RECT 23.18 601.92 933.28 603.63 ;
   RECT 23.18 603.63 933.28 605.34 ;
   RECT 23.18 605.34 933.28 607.05 ;
   RECT 23.18 607.05 933.28 608.76 ;
   RECT 23.18 608.76 933.28 610.47 ;
   RECT 23.18 610.47 933.28 612.18 ;
   RECT 23.18 612.18 933.28 613.89 ;
   RECT 23.18 613.89 933.28 615.6 ;
   RECT 23.18 615.6 933.28 617.31 ;
   RECT 23.18 617.31 933.28 619.02 ;
   RECT 23.18 619.02 933.28 620.73 ;
   RECT 23.18 620.73 933.28 622.44 ;
   RECT 23.18 622.44 933.28 624.15 ;
   RECT 23.18 624.15 933.28 625.86 ;
   RECT 23.18 625.86 933.28 627.57 ;
   RECT 23.18 627.57 933.28 629.28 ;
   RECT 23.18 629.28 933.28 630.99 ;
   RECT 23.18 630.99 933.28 632.7 ;
   RECT 23.18 632.7 933.28 634.41 ;
   RECT 23.18 634.41 933.28 636.12 ;
   RECT 23.18 636.12 933.28 637.83 ;
   RECT 23.18 637.83 933.28 639.54 ;
   RECT 23.18 639.54 933.28 641.25 ;
   RECT 23.18 641.25 933.28 642.96 ;
   RECT 23.18 642.96 933.28 644.67 ;
   RECT 23.18 644.67 933.28 646.38 ;
   RECT 23.18 646.38 933.28 648.09 ;
   RECT 23.18 648.09 933.28 649.8 ;
   RECT 23.18 649.8 933.28 651.51 ;
   RECT 23.18 651.51 933.28 653.22 ;
   RECT 23.18 653.22 933.28 654.93 ;
   RECT 23.18 654.93 933.28 656.64 ;
   RECT 23.18 656.64 933.28 658.35 ;
   RECT 23.18 658.35 933.28 660.06 ;
   RECT 23.18 660.06 933.28 661.77 ;
   RECT 23.18 661.77 933.28 663.48 ;
   RECT 23.18 663.48 933.28 665.19 ;
   RECT 23.18 665.19 933.28 666.9 ;
   RECT 23.18 666.9 933.28 668.61 ;
   RECT 23.18 668.61 933.28 670.32 ;
   RECT 23.18 670.32 933.28 672.03 ;
   RECT 23.18 672.03 933.28 673.74 ;
   RECT 23.18 673.74 933.28 675.45 ;
   RECT 23.18 675.45 933.28 677.16 ;
   RECT 23.18 677.16 933.28 678.87 ;
   RECT 23.18 678.87 933.28 680.58 ;
   RECT 23.18 680.58 933.28 682.29 ;
   RECT 23.18 682.29 933.28 684.0 ;
   RECT 23.18 684.0 933.28 685.71 ;
   RECT 23.18 685.71 933.28 687.42 ;
   RECT 23.18 687.42 933.28 689.13 ;
   RECT 23.18 689.13 933.28 690.84 ;
   RECT 23.18 690.84 933.28 692.55 ;
   RECT 23.18 692.55 933.28 694.26 ;
   RECT 23.18 694.26 933.28 695.97 ;
   RECT 23.18 695.97 933.28 697.68 ;
   RECT 23.18 697.68 933.28 699.39 ;
   RECT 23.18 699.39 933.28 701.1 ;
   RECT 23.18 701.1 933.28 702.81 ;
   RECT 23.18 702.81 933.28 704.52 ;
   RECT 23.18 704.52 933.28 706.23 ;
   RECT 23.18 706.23 933.28 707.94 ;
   RECT 23.18 707.94 933.28 709.65 ;
   RECT 23.18 709.65 933.28 711.36 ;
   RECT 23.18 711.36 933.28 713.07 ;
   RECT 23.18 713.07 933.28 714.78 ;
   RECT 23.18 714.78 933.28 716.49 ;
   RECT 23.18 716.49 933.28 718.2 ;
   RECT 23.18 718.2 933.28 719.91 ;
   RECT 23.18 719.91 933.28 721.62 ;
   RECT 23.18 721.62 933.28 723.33 ;
   RECT 23.18 723.33 933.28 725.04 ;
   RECT 23.18 725.04 933.28 726.75 ;
   RECT 23.18 726.75 933.28 728.46 ;
   RECT 23.18 728.46 933.28 730.17 ;
   RECT 23.18 730.17 933.28 731.88 ;
   RECT 23.18 731.88 933.28 733.59 ;
   RECT 23.18 733.59 933.28 735.3 ;
   RECT 23.18 735.3 933.28 737.01 ;
   RECT 23.18 737.01 933.28 738.72 ;
   RECT 23.18 738.72 933.28 740.43 ;
   RECT 23.18 740.43 933.28 742.14 ;
   RECT 23.18 742.14 933.28 743.85 ;
   RECT 23.18 743.85 933.28 745.56 ;
   RECT 23.18 745.56 933.28 747.27 ;
   RECT 23.18 747.27 933.28 748.98 ;
   RECT 23.18 748.98 933.28 750.69 ;
   RECT 23.18 750.69 933.28 752.4 ;
   RECT 23.18 752.4 933.28 754.11 ;
   RECT 23.18 754.11 933.28 755.82 ;
   RECT 23.18 755.82 933.28 757.53 ;
   RECT 23.18 757.53 933.28 759.24 ;
   RECT 23.18 759.24 933.28 760.95 ;
   RECT 23.18 760.95 933.28 762.66 ;
   RECT 23.18 762.66 933.28 764.37 ;
   RECT 23.18 764.37 933.28 766.08 ;
   RECT 23.18 766.08 933.28 767.79 ;
   RECT 23.18 767.79 933.28 769.5 ;
   RECT 23.18 769.5 933.28 771.21 ;
   RECT 23.18 771.21 933.28 772.92 ;
   RECT 23.18 772.92 933.28 774.63 ;
   RECT 23.18 774.63 933.28 776.34 ;
   RECT 23.18 776.34 933.28 778.05 ;
   RECT 23.18 778.05 933.28 779.76 ;
   RECT 23.18 779.76 933.28 781.47 ;
   RECT 23.18 781.47 933.28 783.18 ;
   RECT 23.18 783.18 933.28 784.89 ;
   RECT 23.18 784.89 933.28 786.6 ;
   RECT 23.18 786.6 933.28 788.31 ;
   RECT 23.18 788.31 933.28 790.02 ;
   RECT 23.18 790.02 933.28 791.73 ;
   RECT 23.18 791.73 933.28 793.44 ;
   RECT 23.18 793.44 933.28 795.15 ;
   RECT 23.18 795.15 933.28 796.86 ;
   RECT 23.18 796.86 933.28 798.57 ;
   RECT 23.18 798.57 933.28 800.28 ;
   RECT 23.18 800.28 933.28 801.99 ;
   RECT 23.18 801.99 933.28 803.7 ;
   RECT 23.18 803.7 933.28 805.41 ;
   RECT 23.18 805.41 933.28 807.12 ;
   RECT 23.18 807.12 933.28 808.83 ;
   RECT 23.18 808.83 933.28 810.54 ;
   RECT 23.18 810.54 933.28 812.25 ;
   RECT 23.18 812.25 933.28 813.96 ;
   RECT 23.18 813.96 933.28 815.67 ;
   RECT 23.18 815.67 933.28 817.38 ;
   RECT 23.18 817.38 933.28 819.09 ;
   RECT 23.18 819.09 933.28 820.8 ;
   RECT 23.18 820.8 933.28 822.51 ;
   RECT 23.18 822.51 933.28 824.22 ;
   RECT 23.18 824.22 933.28 825.93 ;
   RECT 23.18 825.93 933.28 827.64 ;
   RECT 23.18 827.64 933.28 829.35 ;
   RECT 23.18 829.35 933.28 831.06 ;
   RECT 23.18 831.06 933.28 832.77 ;
   RECT 23.18 832.77 933.28 834.48 ;
   RECT 23.18 834.48 933.28 836.19 ;
   RECT 23.18 836.19 933.28 837.9 ;
   RECT 23.18 837.9 933.28 839.61 ;
   RECT 23.18 839.61 933.28 841.32 ;
   RECT 23.18 841.32 933.28 843.03 ;
   RECT 23.18 843.03 933.28 844.74 ;
   RECT 23.18 844.74 933.28 846.45 ;
   RECT 23.18 846.45 933.28 848.16 ;
   RECT 23.18 848.16 933.28 849.87 ;
   RECT 23.18 849.87 933.28 851.58 ;
   RECT 23.18 851.58 933.28 853.29 ;
   RECT 23.18 853.29 933.28 855.0 ;
   RECT 23.18 855.0 933.28 856.71 ;
   RECT 23.18 856.71 933.28 858.42 ;
   RECT 23.18 858.42 933.28 860.13 ;
   RECT 23.18 860.13 933.28 861.84 ;
   RECT 23.18 861.84 933.28 863.55 ;
   RECT 23.18 863.55 933.28 865.26 ;
   RECT 23.18 865.26 933.28 866.97 ;
   RECT 23.18 866.97 933.28 868.68 ;
   RECT 23.18 868.68 933.28 870.39 ;
   RECT 23.18 870.39 933.28 872.1 ;
   RECT 23.18 872.1 933.28 873.81 ;
   RECT 23.18 873.81 933.28 875.52 ;
   RECT 23.18 875.52 933.28 877.23 ;
   RECT 23.18 877.23 933.28 878.94 ;
  LAYER metal4 ;
   RECT 23.18 0.0 933.28 1.71 ;
   RECT 23.18 1.71 933.28 3.42 ;
   RECT 23.18 3.42 933.28 5.13 ;
   RECT 23.18 5.13 933.28 6.84 ;
   RECT 23.18 6.84 933.28 8.55 ;
   RECT 23.18 8.55 933.28 10.26 ;
   RECT 23.18 10.26 933.28 11.97 ;
   RECT 23.18 11.97 933.28 13.68 ;
   RECT 23.18 13.68 933.28 15.39 ;
   RECT 23.18 15.39 933.28 17.1 ;
   RECT 23.18 17.1 933.28 18.81 ;
   RECT 23.18 18.81 933.28 20.52 ;
   RECT 23.18 20.52 933.28 22.23 ;
   RECT 23.18 22.23 933.28 23.94 ;
   RECT 23.18 23.94 933.28 25.65 ;
   RECT 23.18 25.65 933.28 27.36 ;
   RECT 23.18 27.36 933.28 29.07 ;
   RECT 23.18 29.07 933.28 30.78 ;
   RECT 23.18 30.78 933.28 32.49 ;
   RECT 23.18 32.49 933.28 34.2 ;
   RECT 23.18 34.2 933.28 35.91 ;
   RECT 23.18 35.91 933.28 37.62 ;
   RECT 23.18 37.62 933.28 39.33 ;
   RECT 23.18 39.33 933.28 41.04 ;
   RECT 23.18 41.04 933.28 42.75 ;
   RECT 23.18 42.75 933.28 44.46 ;
   RECT 23.18 44.46 933.28 46.17 ;
   RECT 23.18 46.17 933.28 47.88 ;
   RECT 23.18 47.88 933.28 49.59 ;
   RECT 23.18 49.59 933.28 51.3 ;
   RECT 23.18 51.3 933.28 53.01 ;
   RECT 23.18 53.01 933.28 54.72 ;
   RECT 23.18 54.72 933.28 56.43 ;
   RECT 23.18 56.43 933.28 58.14 ;
   RECT 23.18 58.14 933.28 59.85 ;
   RECT 23.18 59.85 933.28 61.56 ;
   RECT 23.18 61.56 933.28 63.27 ;
   RECT 23.18 63.27 933.28 64.98 ;
   RECT 23.18 64.98 933.28 66.69 ;
   RECT 23.18 66.69 933.28 68.4 ;
   RECT 23.18 68.4 933.28 70.11 ;
   RECT 23.18 70.11 933.28 71.82 ;
   RECT 23.18 71.82 933.28 73.53 ;
   RECT 23.18 73.53 933.28 75.24 ;
   RECT 23.18 75.24 933.28 76.95 ;
   RECT 23.18 76.95 933.28 78.66 ;
   RECT 23.18 78.66 933.28 80.37 ;
   RECT 23.18 80.37 933.28 82.08 ;
   RECT 23.18 82.08 933.28 83.79 ;
   RECT 23.18 83.79 933.28 85.5 ;
   RECT 23.18 85.5 933.28 87.21 ;
   RECT 23.18 87.21 933.28 88.92 ;
   RECT 23.18 88.92 933.28 90.63 ;
   RECT 23.18 90.63 933.28 92.34 ;
   RECT 23.18 92.34 933.28 94.05 ;
   RECT 23.18 94.05 933.28 95.76 ;
   RECT 23.18 95.76 933.28 97.47 ;
   RECT 23.18 97.47 933.28 99.18 ;
   RECT 23.18 99.18 933.28 100.89 ;
   RECT 23.18 100.89 933.28 102.6 ;
   RECT 23.18 102.6 933.28 104.31 ;
   RECT 23.18 104.31 933.28 106.02 ;
   RECT 23.18 106.02 933.28 107.73 ;
   RECT 23.18 107.73 933.28 109.44 ;
   RECT 23.18 109.44 933.28 111.15 ;
   RECT 23.18 111.15 933.28 112.86 ;
   RECT 23.18 112.86 933.28 114.57 ;
   RECT 23.18 114.57 933.28 116.28 ;
   RECT 23.18 116.28 933.28 117.99 ;
   RECT 23.18 117.99 933.28 119.7 ;
   RECT 23.18 119.7 933.28 121.41 ;
   RECT 23.18 121.41 933.28 123.12 ;
   RECT 23.18 123.12 933.28 124.83 ;
   RECT 23.18 124.83 933.28 126.54 ;
   RECT 23.18 126.54 933.28 128.25 ;
   RECT 23.18 128.25 933.28 129.96 ;
   RECT 23.18 129.96 933.28 131.67 ;
   RECT 23.18 131.67 933.28 133.38 ;
   RECT 23.18 133.38 933.28 135.09 ;
   RECT 23.18 135.09 933.28 136.8 ;
   RECT 23.18 136.8 933.28 138.51 ;
   RECT 23.18 138.51 933.28 140.22 ;
   RECT 23.18 140.22 933.28 141.93 ;
   RECT 23.18 141.93 933.28 143.64 ;
   RECT 23.18 143.64 933.28 145.35 ;
   RECT 23.18 145.35 933.28 147.06 ;
   RECT 23.18 147.06 933.28 148.77 ;
   RECT 23.18 148.77 933.28 150.48 ;
   RECT 23.18 150.48 933.28 152.19 ;
   RECT 23.18 152.19 933.28 153.9 ;
   RECT 23.18 153.9 933.28 155.61 ;
   RECT 23.18 155.61 933.28 157.32 ;
   RECT 23.18 157.32 933.28 159.03 ;
   RECT 23.18 159.03 933.28 160.74 ;
   RECT 23.18 160.74 933.28 162.45 ;
   RECT 23.18 162.45 933.28 164.16 ;
   RECT 23.18 164.16 933.28 165.87 ;
   RECT 23.18 165.87 933.28 167.58 ;
   RECT 23.18 167.58 933.28 169.29 ;
   RECT 23.18 169.29 933.28 171.0 ;
   RECT 23.18 171.0 933.28 172.71 ;
   RECT 23.18 172.71 933.28 174.42 ;
   RECT 23.18 174.42 933.28 176.13 ;
   RECT 23.18 176.13 933.28 177.84 ;
   RECT 23.18 177.84 933.28 179.55 ;
   RECT 23.18 179.55 933.28 181.26 ;
   RECT 23.18 181.26 933.28 182.97 ;
   RECT 23.18 182.97 933.28 184.68 ;
   RECT 23.18 184.68 933.28 186.39 ;
   RECT 23.18 186.39 933.28 188.1 ;
   RECT 23.18 188.1 933.28 189.81 ;
   RECT 23.18 189.81 933.28 191.52 ;
   RECT 23.18 191.52 933.28 193.23 ;
   RECT 23.18 193.23 933.28 194.94 ;
   RECT 23.18 194.94 933.28 196.65 ;
   RECT 23.18 196.65 933.28 198.36 ;
   RECT 23.18 198.36 933.28 200.07 ;
   RECT 23.18 200.07 933.28 201.78 ;
   RECT 23.18 201.78 933.28 203.49 ;
   RECT 23.18 203.49 933.28 205.2 ;
   RECT 23.18 205.2 933.28 206.91 ;
   RECT 23.18 206.91 933.28 208.62 ;
   RECT 23.18 208.62 933.28 210.33 ;
   RECT 23.18 210.33 933.28 212.04 ;
   RECT 23.18 212.04 933.28 213.75 ;
   RECT 23.18 213.75 933.28 215.46 ;
   RECT 23.18 215.46 933.28 217.17 ;
   RECT 23.18 217.17 933.28 218.88 ;
   RECT 23.18 218.88 933.28 220.59 ;
   RECT 23.18 220.59 933.28 222.3 ;
   RECT 23.18 222.3 933.28 224.01 ;
   RECT 23.18 224.01 933.28 225.72 ;
   RECT 23.18 225.72 933.28 227.43 ;
   RECT 23.18 227.43 933.28 229.14 ;
   RECT 23.18 229.14 933.28 230.85 ;
   RECT 23.18 230.85 933.28 232.56 ;
   RECT 23.18 232.56 933.28 234.27 ;
   RECT 23.18 234.27 933.28 235.98 ;
   RECT 23.18 235.98 933.28 237.69 ;
   RECT 23.18 237.69 933.28 239.4 ;
   RECT 23.18 239.4 933.28 241.11 ;
   RECT 23.18 241.11 933.28 242.82 ;
   RECT 23.18 242.82 933.28 244.53 ;
   RECT 23.18 244.53 933.28 246.24 ;
   RECT 23.18 246.24 933.28 247.95 ;
   RECT 23.18 247.95 933.28 249.66 ;
   RECT 23.18 249.66 933.28 251.37 ;
   RECT 23.18 251.37 933.28 253.08 ;
   RECT 23.18 253.08 933.28 254.79 ;
   RECT 23.18 254.79 933.28 256.5 ;
   RECT 23.18 256.5 933.28 258.21 ;
   RECT 23.18 258.21 933.28 259.92 ;
   RECT 23.18 259.92 933.28 261.63 ;
   RECT 23.18 261.63 933.28 263.34 ;
   RECT 23.18 263.34 933.28 265.05 ;
   RECT 23.18 265.05 933.28 266.76 ;
   RECT 23.18 266.76 933.28 268.47 ;
   RECT 23.18 268.47 933.28 270.18 ;
   RECT 23.18 270.18 933.28 271.89 ;
   RECT 23.18 271.89 933.28 273.6 ;
   RECT 23.18 273.6 933.28 275.31 ;
   RECT 23.18 275.31 933.28 277.02 ;
   RECT 23.18 277.02 933.28 278.73 ;
   RECT 23.18 278.73 933.28 280.44 ;
   RECT 23.18 280.44 933.28 282.15 ;
   RECT 23.18 282.15 933.28 283.86 ;
   RECT 23.18 283.86 933.28 285.57 ;
   RECT 23.18 285.57 933.28 287.28 ;
   RECT 23.18 287.28 933.28 288.99 ;
   RECT 23.18 288.99 933.28 290.7 ;
   RECT 23.18 290.7 933.28 292.41 ;
   RECT 23.18 292.41 933.28 294.12 ;
   RECT 23.18 294.12 933.28 295.83 ;
   RECT 23.18 295.83 933.28 297.54 ;
   RECT 23.18 297.54 933.28 299.25 ;
   RECT 23.18 299.25 933.28 300.96 ;
   RECT 23.18 300.96 933.28 302.67 ;
   RECT 23.18 302.67 933.28 304.38 ;
   RECT 23.18 304.38 933.28 306.09 ;
   RECT 23.18 306.09 933.28 307.8 ;
   RECT 23.18 307.8 933.28 309.51 ;
   RECT 23.18 309.51 933.28 311.22 ;
   RECT 23.18 311.22 933.28 312.93 ;
   RECT 23.18 312.93 933.28 314.64 ;
   RECT 23.18 314.64 933.28 316.35 ;
   RECT 23.18 316.35 933.28 318.06 ;
   RECT 23.18 318.06 933.28 319.77 ;
   RECT 23.18 319.77 933.28 321.48 ;
   RECT 23.18 321.48 933.28 323.19 ;
   RECT 23.18 323.19 933.28 324.9 ;
   RECT 23.18 324.9 933.28 326.61 ;
   RECT 23.18 326.61 933.28 328.32 ;
   RECT 23.18 328.32 933.28 330.03 ;
   RECT 23.18 330.03 933.28 331.74 ;
   RECT 23.18 331.74 933.28 333.45 ;
   RECT 23.18 333.45 933.28 335.16 ;
   RECT 23.18 335.16 933.28 336.87 ;
   RECT 23.18 336.87 933.28 338.58 ;
   RECT 23.18 338.58 933.28 340.29 ;
   RECT 23.18 340.29 933.28 342.0 ;
   RECT 23.18 342.0 933.28 343.71 ;
   RECT 23.18 343.71 933.28 345.42 ;
   RECT 23.18 345.42 933.28 347.13 ;
   RECT 23.18 347.13 933.28 348.84 ;
   RECT 23.18 348.84 933.28 350.55 ;
   RECT 23.18 350.55 933.28 352.26 ;
   RECT 23.18 352.26 933.28 353.97 ;
   RECT 23.18 353.97 933.28 355.68 ;
   RECT 23.18 355.68 933.28 357.39 ;
   RECT 23.18 357.39 933.28 359.1 ;
   RECT 23.18 359.1 933.28 360.81 ;
   RECT 23.18 360.81 933.28 362.52 ;
   RECT 23.18 362.52 933.28 364.23 ;
   RECT 23.18 364.23 933.28 365.94 ;
   RECT 23.18 365.94 933.28 367.65 ;
   RECT 23.18 367.65 933.28 369.36 ;
   RECT 23.18 369.36 933.28 371.07 ;
   RECT 23.18 371.07 933.28 372.78 ;
   RECT 23.18 372.78 933.28 374.49 ;
   RECT 23.18 374.49 933.28 376.2 ;
   RECT 23.18 376.2 933.28 377.91 ;
   RECT 23.18 377.91 933.28 379.62 ;
   RECT 23.18 379.62 933.28 381.33 ;
   RECT 23.18 381.33 933.28 383.04 ;
   RECT 23.18 383.04 933.28 384.75 ;
   RECT 23.18 384.75 933.28 386.46 ;
   RECT 23.18 386.46 933.28 388.17 ;
   RECT 23.18 388.17 933.28 389.88 ;
   RECT 23.18 389.88 933.28 391.59 ;
   RECT 23.18 391.59 933.28 393.3 ;
   RECT 23.18 393.3 933.28 395.01 ;
   RECT 23.18 395.01 933.28 396.72 ;
   RECT 23.18 396.72 933.28 398.43 ;
   RECT 23.18 398.43 933.28 400.14 ;
   RECT 23.18 400.14 933.28 401.85 ;
   RECT 23.18 401.85 933.28 403.56 ;
   RECT 23.18 403.56 933.28 405.27 ;
   RECT 23.18 405.27 933.28 406.98 ;
   RECT 23.18 406.98 933.28 408.69 ;
   RECT 23.18 408.69 933.28 410.4 ;
   RECT 23.18 410.4 933.28 412.11 ;
   RECT 23.18 412.11 933.28 413.82 ;
   RECT 23.18 413.82 933.28 415.53 ;
   RECT 23.18 415.53 933.28 417.24 ;
   RECT 23.18 417.24 933.28 418.95 ;
   RECT 23.18 418.95 933.28 420.66 ;
   RECT 23.18 420.66 933.28 422.37 ;
   RECT 23.18 422.37 933.28 424.08 ;
   RECT 23.18 424.08 933.28 425.79 ;
   RECT 23.18 425.79 933.28 427.5 ;
   RECT 23.18 427.5 933.28 429.21 ;
   RECT 23.18 429.21 933.28 430.92 ;
   RECT 0.0 430.92 933.28 432.63 ;
   RECT 0.0 432.63 933.28 434.34 ;
   RECT 0.0 434.34 933.28 436.05 ;
   RECT 0.0 436.05 933.28 437.76 ;
   RECT 0.0 437.76 933.28 439.47 ;
   RECT 0.0 439.47 933.28 441.18 ;
   RECT 0.0 441.18 933.28 442.89 ;
   RECT 0.0 442.89 933.28 444.6 ;
   RECT 0.0 444.6 933.28 446.31 ;
   RECT 0.0 446.31 933.28 448.02 ;
   RECT 0.0 448.02 933.28 449.73 ;
   RECT 0.0 449.73 933.28 451.44 ;
   RECT 0.0 451.44 933.28 453.15 ;
   RECT 0.0 453.15 933.28 454.86 ;
   RECT 0.0 454.86 933.28 456.57 ;
   RECT 0.0 456.57 933.28 458.28 ;
   RECT 0.0 458.28 933.28 459.99 ;
   RECT 23.18 459.99 933.28 461.7 ;
   RECT 23.18 461.7 933.28 463.41 ;
   RECT 23.18 463.41 933.28 465.12 ;
   RECT 23.18 465.12 933.28 466.83 ;
   RECT 23.18 466.83 933.28 468.54 ;
   RECT 23.18 468.54 933.28 470.25 ;
   RECT 23.18 470.25 933.28 471.96 ;
   RECT 23.18 471.96 933.28 473.67 ;
   RECT 23.18 473.67 933.28 475.38 ;
   RECT 23.18 475.38 933.28 477.09 ;
   RECT 23.18 477.09 933.28 478.8 ;
   RECT 23.18 478.8 933.28 480.51 ;
   RECT 23.18 480.51 933.28 482.22 ;
   RECT 23.18 482.22 933.28 483.93 ;
   RECT 23.18 483.93 933.28 485.64 ;
   RECT 23.18 485.64 933.28 487.35 ;
   RECT 23.18 487.35 933.28 489.06 ;
   RECT 23.18 489.06 933.28 490.77 ;
   RECT 23.18 490.77 933.28 492.48 ;
   RECT 23.18 492.48 933.28 494.19 ;
   RECT 23.18 494.19 933.28 495.9 ;
   RECT 23.18 495.9 933.28 497.61 ;
   RECT 23.18 497.61 933.28 499.32 ;
   RECT 23.18 499.32 933.28 501.03 ;
   RECT 23.18 501.03 933.28 502.74 ;
   RECT 23.18 502.74 933.28 504.45 ;
   RECT 23.18 504.45 933.28 506.16 ;
   RECT 23.18 506.16 933.28 507.87 ;
   RECT 23.18 507.87 933.28 509.58 ;
   RECT 23.18 509.58 933.28 511.29 ;
   RECT 23.18 511.29 933.28 513.0 ;
   RECT 23.18 513.0 933.28 514.71 ;
   RECT 23.18 514.71 933.28 516.42 ;
   RECT 23.18 516.42 933.28 518.13 ;
   RECT 23.18 518.13 933.28 519.84 ;
   RECT 23.18 519.84 933.28 521.55 ;
   RECT 23.18 521.55 933.28 523.26 ;
   RECT 23.18 523.26 933.28 524.97 ;
   RECT 23.18 524.97 933.28 526.68 ;
   RECT 23.18 526.68 933.28 528.39 ;
   RECT 23.18 528.39 933.28 530.1 ;
   RECT 23.18 530.1 933.28 531.81 ;
   RECT 23.18 531.81 933.28 533.52 ;
   RECT 23.18 533.52 933.28 535.23 ;
   RECT 23.18 535.23 933.28 536.94 ;
   RECT 23.18 536.94 933.28 538.65 ;
   RECT 23.18 538.65 933.28 540.36 ;
   RECT 23.18 540.36 933.28 542.07 ;
   RECT 23.18 542.07 933.28 543.78 ;
   RECT 23.18 543.78 933.28 545.49 ;
   RECT 23.18 545.49 933.28 547.2 ;
   RECT 23.18 547.2 933.28 548.91 ;
   RECT 23.18 548.91 933.28 550.62 ;
   RECT 23.18 550.62 933.28 552.33 ;
   RECT 23.18 552.33 933.28 554.04 ;
   RECT 23.18 554.04 933.28 555.75 ;
   RECT 23.18 555.75 933.28 557.46 ;
   RECT 23.18 557.46 933.28 559.17 ;
   RECT 23.18 559.17 933.28 560.88 ;
   RECT 23.18 560.88 933.28 562.59 ;
   RECT 23.18 562.59 933.28 564.3 ;
   RECT 23.18 564.3 933.28 566.01 ;
   RECT 23.18 566.01 933.28 567.72 ;
   RECT 23.18 567.72 933.28 569.43 ;
   RECT 23.18 569.43 933.28 571.14 ;
   RECT 23.18 571.14 933.28 572.85 ;
   RECT 23.18 572.85 933.28 574.56 ;
   RECT 23.18 574.56 933.28 576.27 ;
   RECT 23.18 576.27 933.28 577.98 ;
   RECT 23.18 577.98 933.28 579.69 ;
   RECT 23.18 579.69 933.28 581.4 ;
   RECT 23.18 581.4 933.28 583.11 ;
   RECT 23.18 583.11 933.28 584.82 ;
   RECT 23.18 584.82 933.28 586.53 ;
   RECT 23.18 586.53 933.28 588.24 ;
   RECT 23.18 588.24 933.28 589.95 ;
   RECT 23.18 589.95 933.28 591.66 ;
   RECT 23.18 591.66 933.28 593.37 ;
   RECT 23.18 593.37 933.28 595.08 ;
   RECT 23.18 595.08 933.28 596.79 ;
   RECT 23.18 596.79 933.28 598.5 ;
   RECT 23.18 598.5 933.28 600.21 ;
   RECT 23.18 600.21 933.28 601.92 ;
   RECT 23.18 601.92 933.28 603.63 ;
   RECT 23.18 603.63 933.28 605.34 ;
   RECT 23.18 605.34 933.28 607.05 ;
   RECT 23.18 607.05 933.28 608.76 ;
   RECT 23.18 608.76 933.28 610.47 ;
   RECT 23.18 610.47 933.28 612.18 ;
   RECT 23.18 612.18 933.28 613.89 ;
   RECT 23.18 613.89 933.28 615.6 ;
   RECT 23.18 615.6 933.28 617.31 ;
   RECT 23.18 617.31 933.28 619.02 ;
   RECT 23.18 619.02 933.28 620.73 ;
   RECT 23.18 620.73 933.28 622.44 ;
   RECT 23.18 622.44 933.28 624.15 ;
   RECT 23.18 624.15 933.28 625.86 ;
   RECT 23.18 625.86 933.28 627.57 ;
   RECT 23.18 627.57 933.28 629.28 ;
   RECT 23.18 629.28 933.28 630.99 ;
   RECT 23.18 630.99 933.28 632.7 ;
   RECT 23.18 632.7 933.28 634.41 ;
   RECT 23.18 634.41 933.28 636.12 ;
   RECT 23.18 636.12 933.28 637.83 ;
   RECT 23.18 637.83 933.28 639.54 ;
   RECT 23.18 639.54 933.28 641.25 ;
   RECT 23.18 641.25 933.28 642.96 ;
   RECT 23.18 642.96 933.28 644.67 ;
   RECT 23.18 644.67 933.28 646.38 ;
   RECT 23.18 646.38 933.28 648.09 ;
   RECT 23.18 648.09 933.28 649.8 ;
   RECT 23.18 649.8 933.28 651.51 ;
   RECT 23.18 651.51 933.28 653.22 ;
   RECT 23.18 653.22 933.28 654.93 ;
   RECT 23.18 654.93 933.28 656.64 ;
   RECT 23.18 656.64 933.28 658.35 ;
   RECT 23.18 658.35 933.28 660.06 ;
   RECT 23.18 660.06 933.28 661.77 ;
   RECT 23.18 661.77 933.28 663.48 ;
   RECT 23.18 663.48 933.28 665.19 ;
   RECT 23.18 665.19 933.28 666.9 ;
   RECT 23.18 666.9 933.28 668.61 ;
   RECT 23.18 668.61 933.28 670.32 ;
   RECT 23.18 670.32 933.28 672.03 ;
   RECT 23.18 672.03 933.28 673.74 ;
   RECT 23.18 673.74 933.28 675.45 ;
   RECT 23.18 675.45 933.28 677.16 ;
   RECT 23.18 677.16 933.28 678.87 ;
   RECT 23.18 678.87 933.28 680.58 ;
   RECT 23.18 680.58 933.28 682.29 ;
   RECT 23.18 682.29 933.28 684.0 ;
   RECT 23.18 684.0 933.28 685.71 ;
   RECT 23.18 685.71 933.28 687.42 ;
   RECT 23.18 687.42 933.28 689.13 ;
   RECT 23.18 689.13 933.28 690.84 ;
   RECT 23.18 690.84 933.28 692.55 ;
   RECT 23.18 692.55 933.28 694.26 ;
   RECT 23.18 694.26 933.28 695.97 ;
   RECT 23.18 695.97 933.28 697.68 ;
   RECT 23.18 697.68 933.28 699.39 ;
   RECT 23.18 699.39 933.28 701.1 ;
   RECT 23.18 701.1 933.28 702.81 ;
   RECT 23.18 702.81 933.28 704.52 ;
   RECT 23.18 704.52 933.28 706.23 ;
   RECT 23.18 706.23 933.28 707.94 ;
   RECT 23.18 707.94 933.28 709.65 ;
   RECT 23.18 709.65 933.28 711.36 ;
   RECT 23.18 711.36 933.28 713.07 ;
   RECT 23.18 713.07 933.28 714.78 ;
   RECT 23.18 714.78 933.28 716.49 ;
   RECT 23.18 716.49 933.28 718.2 ;
   RECT 23.18 718.2 933.28 719.91 ;
   RECT 23.18 719.91 933.28 721.62 ;
   RECT 23.18 721.62 933.28 723.33 ;
   RECT 23.18 723.33 933.28 725.04 ;
   RECT 23.18 725.04 933.28 726.75 ;
   RECT 23.18 726.75 933.28 728.46 ;
   RECT 23.18 728.46 933.28 730.17 ;
   RECT 23.18 730.17 933.28 731.88 ;
   RECT 23.18 731.88 933.28 733.59 ;
   RECT 23.18 733.59 933.28 735.3 ;
   RECT 23.18 735.3 933.28 737.01 ;
   RECT 23.18 737.01 933.28 738.72 ;
   RECT 23.18 738.72 933.28 740.43 ;
   RECT 23.18 740.43 933.28 742.14 ;
   RECT 23.18 742.14 933.28 743.85 ;
   RECT 23.18 743.85 933.28 745.56 ;
   RECT 23.18 745.56 933.28 747.27 ;
   RECT 23.18 747.27 933.28 748.98 ;
   RECT 23.18 748.98 933.28 750.69 ;
   RECT 23.18 750.69 933.28 752.4 ;
   RECT 23.18 752.4 933.28 754.11 ;
   RECT 23.18 754.11 933.28 755.82 ;
   RECT 23.18 755.82 933.28 757.53 ;
   RECT 23.18 757.53 933.28 759.24 ;
   RECT 23.18 759.24 933.28 760.95 ;
   RECT 23.18 760.95 933.28 762.66 ;
   RECT 23.18 762.66 933.28 764.37 ;
   RECT 23.18 764.37 933.28 766.08 ;
   RECT 23.18 766.08 933.28 767.79 ;
   RECT 23.18 767.79 933.28 769.5 ;
   RECT 23.18 769.5 933.28 771.21 ;
   RECT 23.18 771.21 933.28 772.92 ;
   RECT 23.18 772.92 933.28 774.63 ;
   RECT 23.18 774.63 933.28 776.34 ;
   RECT 23.18 776.34 933.28 778.05 ;
   RECT 23.18 778.05 933.28 779.76 ;
   RECT 23.18 779.76 933.28 781.47 ;
   RECT 23.18 781.47 933.28 783.18 ;
   RECT 23.18 783.18 933.28 784.89 ;
   RECT 23.18 784.89 933.28 786.6 ;
   RECT 23.18 786.6 933.28 788.31 ;
   RECT 23.18 788.31 933.28 790.02 ;
   RECT 23.18 790.02 933.28 791.73 ;
   RECT 23.18 791.73 933.28 793.44 ;
   RECT 23.18 793.44 933.28 795.15 ;
   RECT 23.18 795.15 933.28 796.86 ;
   RECT 23.18 796.86 933.28 798.57 ;
   RECT 23.18 798.57 933.28 800.28 ;
   RECT 23.18 800.28 933.28 801.99 ;
   RECT 23.18 801.99 933.28 803.7 ;
   RECT 23.18 803.7 933.28 805.41 ;
   RECT 23.18 805.41 933.28 807.12 ;
   RECT 23.18 807.12 933.28 808.83 ;
   RECT 23.18 808.83 933.28 810.54 ;
   RECT 23.18 810.54 933.28 812.25 ;
   RECT 23.18 812.25 933.28 813.96 ;
   RECT 23.18 813.96 933.28 815.67 ;
   RECT 23.18 815.67 933.28 817.38 ;
   RECT 23.18 817.38 933.28 819.09 ;
   RECT 23.18 819.09 933.28 820.8 ;
   RECT 23.18 820.8 933.28 822.51 ;
   RECT 23.18 822.51 933.28 824.22 ;
   RECT 23.18 824.22 933.28 825.93 ;
   RECT 23.18 825.93 933.28 827.64 ;
   RECT 23.18 827.64 933.28 829.35 ;
   RECT 23.18 829.35 933.28 831.06 ;
   RECT 23.18 831.06 933.28 832.77 ;
   RECT 23.18 832.77 933.28 834.48 ;
   RECT 23.18 834.48 933.28 836.19 ;
   RECT 23.18 836.19 933.28 837.9 ;
   RECT 23.18 837.9 933.28 839.61 ;
   RECT 23.18 839.61 933.28 841.32 ;
   RECT 23.18 841.32 933.28 843.03 ;
   RECT 23.18 843.03 933.28 844.74 ;
   RECT 23.18 844.74 933.28 846.45 ;
   RECT 23.18 846.45 933.28 848.16 ;
   RECT 23.18 848.16 933.28 849.87 ;
   RECT 23.18 849.87 933.28 851.58 ;
   RECT 23.18 851.58 933.28 853.29 ;
   RECT 23.18 853.29 933.28 855.0 ;
   RECT 23.18 855.0 933.28 856.71 ;
   RECT 23.18 856.71 933.28 858.42 ;
   RECT 23.18 858.42 933.28 860.13 ;
   RECT 23.18 860.13 933.28 861.84 ;
   RECT 23.18 861.84 933.28 863.55 ;
   RECT 23.18 863.55 933.28 865.26 ;
   RECT 23.18 865.26 933.28 866.97 ;
   RECT 23.18 866.97 933.28 868.68 ;
   RECT 23.18 868.68 933.28 870.39 ;
   RECT 23.18 870.39 933.28 872.1 ;
   RECT 23.18 872.1 933.28 873.81 ;
   RECT 23.18 873.81 933.28 875.52 ;
   RECT 23.18 875.52 933.28 877.23 ;
   RECT 23.18 877.23 933.28 878.94 ;
 END
END block_2456x4626_834

MACRO block_416x441_112
 CLASS BLOCK ;
 FOREIGN block_416x441_112 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 158.08 BY 83.79 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 64.315 154.945 64.885 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 20.615 154.945 21.185 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 4.655 3.325 5.225 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 6.175 3.325 6.745 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 7.315 3.325 7.885 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 8.075 3.325 8.645 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 9.215 3.325 9.785 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 10.735 3.325 11.305 ;
  END
 END o7
 PIN o8
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 11.875 3.325 12.445 ;
  END
 END o8
 PIN o9
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 12.635 3.325 13.205 ;
  END
 END o9
 PIN o10
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 24.415 3.325 24.985 ;
  END
 END o10
 PIN o11
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 25.555 3.325 26.125 ;
  END
 END o11
 PIN o12
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 26.315 3.325 26.885 ;
  END
 END o12
 PIN o13
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 27.455 3.325 28.025 ;
  END
 END o13
 PIN o14
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 28.975 3.325 29.545 ;
  END
 END o14
 PIN o15
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 22.895 3.325 23.465 ;
  END
 END o15
 PIN o16
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 32.015 3.325 32.585 ;
  END
 END o16
 PIN o17
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 33.535 3.325 34.105 ;
  END
 END o17
 PIN o18
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 34.295 3.325 34.865 ;
  END
 END o18
 PIN o19
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 35.055 3.325 35.625 ;
  END
 END o19
 PIN o20
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 35.815 3.325 36.385 ;
  END
 END o20
 PIN o21
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 30.875 3.325 31.445 ;
  END
 END o21
 PIN o22
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 38.855 3.325 39.425 ;
  END
 END o22
 PIN o23
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 39.615 3.325 40.185 ;
  END
 END o23
 PIN o24
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 40.375 3.325 40.945 ;
  END
 END o24
 PIN o25
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 41.135 3.325 41.705 ;
  END
 END o25
 PIN o26
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 42.655 3.325 43.225 ;
  END
 END o26
 PIN o27
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 38.095 3.325 38.665 ;
  END
 END o27
 PIN o28
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 44.935 3.325 45.505 ;
  END
 END o28
 PIN o29
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 45.695 3.325 46.265 ;
  END
 END o29
 PIN o30
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 47.215 3.325 47.785 ;
  END
 END o30
 PIN o31
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 47.975 3.325 48.545 ;
  END
 END o31
 PIN o32
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 48.735 3.325 49.305 ;
  END
 END o32
 PIN o33
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 44.175 3.325 44.745 ;
  END
 END o33
 PIN o34
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 51.775 3.325 52.345 ;
  END
 END o34
 PIN o35
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 52.535 3.325 53.105 ;
  END
 END o35
 PIN o36
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 53.295 3.325 53.865 ;
  END
 END o36
 PIN o37
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 54.055 3.325 54.625 ;
  END
 END o37
 PIN o38
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 54.815 3.325 55.385 ;
  END
 END o38
 PIN o39
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 50.255 3.325 50.825 ;
  END
 END o39
 PIN o40
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 57.855 3.325 58.425 ;
  END
 END o40
 PIN o41
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 58.615 3.325 59.185 ;
  END
 END o41
 PIN o42
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 59.375 3.325 59.945 ;
  END
 END o42
 PIN o43
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 60.895 3.325 61.465 ;
  END
 END o43
 PIN o44
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 61.655 3.325 62.225 ;
  END
 END o44
 PIN o45
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 57.095 3.325 57.665 ;
  END
 END o45
 PIN o46
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 63.935 3.325 64.505 ;
  END
 END o46
 PIN o47
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 65.455 3.325 66.025 ;
  END
 END o47
 PIN o48
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 66.215 3.325 66.785 ;
  END
 END o48
 PIN o49
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 66.975 3.325 67.545 ;
  END
 END o49
 PIN o50
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 67.735 3.325 68.305 ;
  END
 END o50
 PIN o51
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 63.175 3.325 63.745 ;
  END
 END o51
 PIN o52
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 70.775 3.325 71.345 ;
  END
 END o52
 PIN o53
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 71.535 3.325 72.105 ;
  END
 END o53
 PIN o54
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 72.295 3.325 72.865 ;
  END
 END o54
 PIN o55
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 72.675 4.085 73.245 ;
  END
 END o55
 PIN o56
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 73.055 3.325 73.625 ;
  END
 END o56
 PIN o57
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 70.015 3.325 70.585 ;
  END
 END o57
 PIN o58
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 24.415 154.945 24.985 ;
  END
 END o58
 PIN o59
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 25.175 154.945 25.745 ;
  END
 END o59
 PIN o60
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 25.935 154.945 26.505 ;
  END
 END o60
 PIN o61
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 26.695 154.945 27.265 ;
  END
 END o61
 PIN o62
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 27.455 154.945 28.025 ;
  END
 END o62
 PIN o63
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 22.895 154.945 23.465 ;
  END
 END o63
 PIN o64
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 29.735 154.945 30.305 ;
  END
 END o64
 PIN o65
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 30.495 154.945 31.065 ;
  END
 END o65
 PIN o66
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 31.255 154.945 31.825 ;
  END
 END o66
 PIN o67
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 32.015 154.945 32.585 ;
  END
 END o67
 PIN o68
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 33.535 154.945 34.105 ;
  END
 END o68
 PIN o69
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 28.975 154.945 29.545 ;
  END
 END o69
 PIN o70
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 22.135 154.945 22.705 ;
  END
 END o70
 PIN o71
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 74.955 3.325 75.525 ;
  END
 END o71
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 51.775 154.945 52.345 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 66.975 154.945 67.545 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 49.495 154.945 50.065 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 50.255 154.945 50.825 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 54.055 154.945 54.625 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 53.295 154.945 53.865 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 47.215 154.945 47.785 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 47.975 154.945 48.545 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 21.375 154.945 21.945 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 74.575 4.085 75.145 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 57.095 154.945 57.665 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 57.855 154.945 58.425 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 58.615 154.945 59.185 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 59.375 154.945 59.945 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 60.895 154.945 61.465 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 61.655 154.945 62.225 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 62.415 154.945 62.985 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 63.175 154.945 63.745 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 3.135 154.945 3.705 ;
  END
 END i18
 PIN i19
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 3.895 154.945 4.465 ;
  END
 END i19
 PIN i20
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 4.655 154.945 5.225 ;
  END
 END i20
 PIN i21
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 6.175 154.945 6.745 ;
  END
 END i21
 PIN i22
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 6.935 154.945 7.505 ;
  END
 END i22
 PIN i23
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 7.695 154.945 8.265 ;
  END
 END i23
 PIN i24
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 3.515 3.325 4.085 ;
  END
 END i24
 PIN i25
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 19.855 154.945 20.425 ;
  END
 END i25
 PIN i26
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 18.335 154.945 18.905 ;
  END
 END i26
 PIN i27
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 17.575 154.945 18.145 ;
  END
 END i27
 PIN i28
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 48.735 154.945 49.305 ;
  END
 END i28
 PIN i29
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 45.695 154.945 46.265 ;
  END
 END i29
 PIN i30
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 44.935 154.945 45.505 ;
  END
 END i30
 PIN i31
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 8.455 154.945 9.025 ;
  END
 END i31
 PIN i32
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 9.215 154.945 9.785 ;
  END
 END i32
 PIN i33
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 10.735 154.945 11.305 ;
  END
 END i33
 PIN i34
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 11.495 154.945 12.065 ;
  END
 END i34
 PIN i35
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 12.255 154.945 12.825 ;
  END
 END i35
 PIN i36
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 13.015 154.945 13.585 ;
  END
 END i36
 PIN i37
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 13.775 154.945 14.345 ;
  END
 END i37
 PIN i38
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 15.295 154.945 15.865 ;
  END
 END i38
 PIN i39
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 16.055 154.945 16.625 ;
  END
 END i39
 OBS
  LAYER metal1 ;
   RECT 0 0 158.08 83.79 ;
  LAYER via1 ;
   RECT 0 0 158.08 83.79 ;
  LAYER metal2 ;
   RECT 0 0 158.08 83.79 ;
  LAYER via2 ;
   RECT 0 0 158.08 83.79 ;
  LAYER metal3 ;
   RECT 0 0 158.08 83.79 ;
  LAYER via3 ;
   RECT 0 0 158.08 83.79 ;
  LAYER metal4 ;
   RECT 0 0 158.08 83.79 ;
 END
END block_416x441_112

MACRO block_126x351_27
 CLASS BLOCK ;
 FOREIGN block_126x351_27 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 47.88 BY 66.69 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 2.565 9.785 3.135 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 8.265 9.785 8.835 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 14.155 9.785 14.725 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 19.855 9.785 20.425 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 57.095 9.785 57.665 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 62.795 9.785 63.365 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 51.395 9.785 51.965 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 46.075 1.045 46.645 1.615 ;
  END
 END o7
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 46.075 27.645 46.645 28.215 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 46.075 28.975 46.645 29.545 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 39.995 27.835 40.565 28.405 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 46.075 36.955 46.645 37.525 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 28.405 9.785 28.975 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 46.075 44.365 46.645 44.935 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 46.075 34.485 46.645 35.055 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 46.075 35.625 46.645 36.195 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 35.435 9.785 36.005 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 8.455 42.275 9.025 42.845 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 39.235 9.785 39.805 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 45.315 37.525 45.885 38.095 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 46.075 62.415 46.645 62.985 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 46.075 56.715 46.645 57.285 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 46.075 51.015 46.645 51.585 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 46.075 20.235 46.645 20.805 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 46.075 14.535 46.645 15.105 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 46.075 8.835 46.645 9.405 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 46.075 2.945 46.645 3.515 ;
  END
 END i18
 OBS
  LAYER metal1 ;
   RECT 0 0 47.88 66.69 ;
  LAYER via1 ;
   RECT 0 0 47.88 66.69 ;
  LAYER metal2 ;
   RECT 0 0 47.88 66.69 ;
  LAYER via2 ;
   RECT 0 0 47.88 66.69 ;
  LAYER metal3 ;
   RECT 0 0 47.88 66.69 ;
  LAYER via3 ;
   RECT 0 0 47.88 66.69 ;
  LAYER metal4 ;
   RECT 0 0 47.88 66.69 ;
 END
END block_126x351_27

MACRO block_533x1539_269
 CLASS BLOCK ;
 FOREIGN block_533x1539_269 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 202.54 BY 292.41 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 4.275 26.885 4.845 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 8.455 26.885 9.025 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 45.125 26.885 45.695 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 49.305 26.885 49.875 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 53.295 26.885 53.865 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 57.475 26.885 58.045 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 79.705 26.885 80.275 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 83.885 26.885 84.455 ;
  END
 END o7
 PIN o8
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 87.875 26.885 88.445 ;
  END
 END o8
 PIN o9
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 92.055 26.885 92.625 ;
  END
 END o9
 PIN o10
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 96.045 26.885 96.615 ;
  END
 END o10
 PIN o11
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 100.225 26.885 100.795 ;
  END
 END o11
 PIN o12
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 12.445 26.885 13.015 ;
  END
 END o12
 PIN o13
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 104.215 26.885 104.785 ;
  END
 END o13
 PIN o14
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 108.395 26.885 108.965 ;
  END
 END o14
 PIN o15
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 112.385 26.885 112.955 ;
  END
 END o15
 PIN o16
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 116.565 26.885 117.135 ;
  END
 END o16
 PIN o17
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 120.555 26.885 121.125 ;
  END
 END o17
 PIN o18
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 124.735 26.885 125.305 ;
  END
 END o18
 PIN o19
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 128.725 26.885 129.295 ;
  END
 END o19
 PIN o20
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 132.905 26.885 133.475 ;
  END
 END o20
 PIN o21
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 161.025 26.885 161.595 ;
  END
 END o21
 PIN o22
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 165.205 26.885 165.775 ;
  END
 END o22
 PIN o23
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 16.625 26.885 17.195 ;
  END
 END o23
 PIN o24
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 169.195 26.885 169.765 ;
  END
 END o24
 PIN o25
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 173.375 26.885 173.945 ;
  END
 END o25
 PIN o26
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 177.365 26.885 177.935 ;
  END
 END o26
 PIN o27
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 181.545 26.885 182.115 ;
  END
 END o27
 PIN o28
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 185.535 26.885 186.105 ;
  END
 END o28
 PIN o29
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 189.715 26.885 190.285 ;
  END
 END o29
 PIN o30
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 193.705 26.885 194.275 ;
  END
 END o30
 PIN o31
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 197.885 26.885 198.455 ;
  END
 END o31
 PIN o32
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 201.875 26.885 202.445 ;
  END
 END o32
 PIN o33
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 206.055 26.885 206.625 ;
  END
 END o33
 PIN o34
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 20.615 26.885 21.185 ;
  END
 END o34
 PIN o35
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 210.045 26.885 210.615 ;
  END
 END o35
 PIN o36
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 214.225 26.885 214.795 ;
  END
 END o36
 PIN o37
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 236.455 26.885 237.025 ;
  END
 END o37
 PIN o38
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 240.635 26.885 241.205 ;
  END
 END o38
 PIN o39
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 244.625 26.885 245.195 ;
  END
 END o39
 PIN o40
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 248.805 26.885 249.375 ;
  END
 END o40
 PIN o41
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 252.795 26.885 253.365 ;
  END
 END o41
 PIN o42
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 256.975 26.885 257.545 ;
  END
 END o42
 PIN o43
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 260.965 26.885 261.535 ;
  END
 END o43
 PIN o44
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 265.145 26.885 265.715 ;
  END
 END o44
 PIN o45
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 24.795 26.885 25.365 ;
  END
 END o45
 PIN o46
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 269.135 26.885 269.705 ;
  END
 END o46
 PIN o47
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 273.315 26.885 273.885 ;
  END
 END o47
 PIN o48
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 277.305 26.885 277.875 ;
  END
 END o48
 PIN o49
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 281.485 26.885 282.055 ;
  END
 END o49
 PIN o50
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 285.475 26.885 286.045 ;
  END
 END o50
 PIN o51
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 28.785 26.885 29.355 ;
  END
 END o51
 PIN o52
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 32.965 26.885 33.535 ;
  END
 END o52
 PIN o53
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 36.955 26.885 37.525 ;
  END
 END o53
 PIN o54
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 41.135 26.885 41.705 ;
  END
 END o54
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 135.755 3.705 136.325 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 152.855 3.705 153.425 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 141.075 3.705 141.645 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 136.135 4.465 136.705 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 135.375 4.465 135.945 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 134.995 3.705 135.565 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 144.685 3.705 145.255 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 157.795 3.705 158.365 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 152.475 4.465 153.045 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 152.095 3.705 152.665 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 154.185 3.705 154.755 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 156.655 3.705 157.225 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 158.175 4.465 158.745 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 13.015 134.615 13.585 135.185 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 13.015 147.915 13.585 148.485 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 2.565 26.885 3.135 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 6.745 26.885 7.315 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 43.415 26.885 43.985 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 47.595 26.885 48.165 ;
  END
 END i18
 PIN i19
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 51.585 26.885 52.155 ;
  END
 END i19
 PIN i20
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 55.765 26.885 56.335 ;
  END
 END i20
 PIN i21
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 77.995 26.885 78.565 ;
  END
 END i21
 PIN i22
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 82.175 26.885 82.745 ;
  END
 END i22
 PIN i23
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 86.165 26.885 86.735 ;
  END
 END i23
 PIN i24
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 90.345 26.885 90.915 ;
  END
 END i24
 PIN i25
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 94.335 26.885 94.905 ;
  END
 END i25
 PIN i26
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 98.515 26.885 99.085 ;
  END
 END i26
 PIN i27
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 10.735 26.885 11.305 ;
  END
 END i27
 PIN i28
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 102.505 26.885 103.075 ;
  END
 END i28
 PIN i29
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 106.685 26.885 107.255 ;
  END
 END i29
 PIN i30
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 110.675 26.885 111.245 ;
  END
 END i30
 PIN i31
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 114.855 26.885 115.425 ;
  END
 END i31
 PIN i32
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 118.845 26.885 119.415 ;
  END
 END i32
 PIN i33
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 123.025 26.885 123.595 ;
  END
 END i33
 PIN i34
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 127.015 26.885 127.585 ;
  END
 END i34
 PIN i35
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 131.195 26.885 131.765 ;
  END
 END i35
 PIN i36
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 162.735 26.885 163.305 ;
  END
 END i36
 PIN i37
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 166.915 26.885 167.485 ;
  END
 END i37
 PIN i38
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 14.915 26.885 15.485 ;
  END
 END i38
 PIN i39
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 170.905 26.885 171.475 ;
  END
 END i39
 PIN i40
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 175.085 26.885 175.655 ;
  END
 END i40
 PIN i41
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 179.075 26.885 179.645 ;
  END
 END i41
 PIN i42
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 183.255 26.885 183.825 ;
  END
 END i42
 PIN i43
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 187.245 26.885 187.815 ;
  END
 END i43
 PIN i44
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 191.425 26.885 191.995 ;
  END
 END i44
 PIN i45
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 195.415 26.885 195.985 ;
  END
 END i45
 PIN i46
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 199.595 26.885 200.165 ;
  END
 END i46
 PIN i47
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 203.585 26.885 204.155 ;
  END
 END i47
 PIN i48
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 207.765 26.885 208.335 ;
  END
 END i48
 PIN i49
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 18.905 26.885 19.475 ;
  END
 END i49
 PIN i50
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 211.755 26.885 212.325 ;
  END
 END i50
 PIN i51
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 215.935 26.885 216.505 ;
  END
 END i51
 PIN i52
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 238.165 26.885 238.735 ;
  END
 END i52
 PIN i53
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 242.345 26.885 242.915 ;
  END
 END i53
 PIN i54
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 246.335 26.885 246.905 ;
  END
 END i54
 PIN i55
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 250.515 26.885 251.085 ;
  END
 END i55
 PIN i56
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 254.505 26.885 255.075 ;
  END
 END i56
 PIN i57
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 258.685 26.885 259.255 ;
  END
 END i57
 PIN i58
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 262.675 26.885 263.245 ;
  END
 END i58
 PIN i59
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 266.855 26.885 267.425 ;
  END
 END i59
 PIN i60
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 23.085 26.885 23.655 ;
  END
 END i60
 PIN i61
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 270.845 26.885 271.415 ;
  END
 END i61
 PIN i62
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 275.025 26.885 275.595 ;
  END
 END i62
 PIN i63
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 279.015 26.885 279.585 ;
  END
 END i63
 PIN i64
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 283.195 26.885 283.765 ;
  END
 END i64
 PIN i65
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 287.185 26.885 287.755 ;
  END
 END i65
 PIN i66
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 27.075 26.885 27.645 ;
  END
 END i66
 PIN i67
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 31.255 26.885 31.825 ;
  END
 END i67
 PIN i68
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 35.245 26.885 35.815 ;
  END
 END i68
 PIN i69
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 39.425 26.885 39.995 ;
  END
 END i69
 PIN i70
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 33.535 27.645 34.105 ;
  END
 END i70
 PIN i71
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 37.525 27.645 38.095 ;
  END
 END i71
 PIN i72
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 41.705 27.645 42.275 ;
  END
 END i72
 PIN i73
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 25.365 27.645 25.935 ;
  END
 END i73
 PIN i74
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 100.795 27.645 101.365 ;
  END
 END i74
 PIN i75
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 104.785 27.645 105.355 ;
  END
 END i75
 PIN i76
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 108.965 27.645 109.535 ;
  END
 END i76
 PIN i77
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 112.955 27.645 113.525 ;
  END
 END i77
 PIN i78
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 193.135 27.645 193.705 ;
  END
 END i78
 PIN i79
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 189.145 27.645 189.715 ;
  END
 END i79
 PIN i80
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 184.965 27.645 185.535 ;
  END
 END i80
 PIN i81
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 180.975 27.645 181.545 ;
  END
 END i81
 PIN i82
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 260.395 27.645 260.965 ;
  END
 END i82
 PIN i83
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 256.405 27.645 256.975 ;
  END
 END i83
 PIN i84
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 252.225 27.645 252.795 ;
  END
 END i84
 PIN i85
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 268.565 27.645 269.135 ;
  END
 END i85
 PIN i86
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 29.355 27.645 29.925 ;
  END
 END i86
 PIN i87
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 96.615 27.645 97.185 ;
  END
 END i87
 PIN i88
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 197.315 27.645 197.885 ;
  END
 END i88
 PIN i89
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 264.575 27.645 265.145 ;
  END
 END i89
 PIN i90
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 17.955 134.615 18.525 135.185 ;
  END
 END i90
 PIN i91
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 17.955 147.915 18.525 148.485 ;
  END
 END i91
 PIN i92
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 3.135 27.645 3.705 ;
  END
 END i92
 PIN i93
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 7.315 27.645 7.885 ;
  END
 END i93
 PIN i94
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 43.985 27.645 44.555 ;
  END
 END i94
 PIN i95
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 48.165 27.645 48.735 ;
  END
 END i95
 PIN i96
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 52.155 27.645 52.725 ;
  END
 END i96
 PIN i97
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 56.335 27.645 56.905 ;
  END
 END i97
 PIN i98
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 78.565 27.645 79.135 ;
  END
 END i98
 PIN i99
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 82.745 27.645 83.315 ;
  END
 END i99
 PIN i100
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 86.735 27.645 87.305 ;
  END
 END i100
 PIN i101
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 90.915 27.645 91.485 ;
  END
 END i101
 PIN i102
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 94.905 27.645 95.475 ;
  END
 END i102
 PIN i103
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 99.085 27.645 99.655 ;
  END
 END i103
 PIN i104
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 11.305 27.645 11.875 ;
  END
 END i104
 PIN i105
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 103.075 27.645 103.645 ;
  END
 END i105
 PIN i106
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 107.255 27.645 107.825 ;
  END
 END i106
 PIN i107
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 111.245 27.645 111.815 ;
  END
 END i107
 PIN i108
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 115.425 27.645 115.995 ;
  END
 END i108
 PIN i109
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 119.415 27.645 119.985 ;
  END
 END i109
 PIN i110
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 123.595 27.645 124.165 ;
  END
 END i110
 PIN i111
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 127.585 27.645 128.155 ;
  END
 END i111
 PIN i112
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 131.765 27.645 132.335 ;
  END
 END i112
 PIN i113
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 162.165 27.645 162.735 ;
  END
 END i113
 PIN i114
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 166.345 27.645 166.915 ;
  END
 END i114
 PIN i115
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 15.485 27.645 16.055 ;
  END
 END i115
 PIN i116
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 170.335 27.645 170.905 ;
  END
 END i116
 PIN i117
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 174.515 27.645 175.085 ;
  END
 END i117
 PIN i118
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 178.505 27.645 179.075 ;
  END
 END i118
 PIN i119
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 182.685 27.645 183.255 ;
  END
 END i119
 PIN i120
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 186.675 27.645 187.245 ;
  END
 END i120
 PIN i121
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 190.855 27.645 191.425 ;
  END
 END i121
 PIN i122
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 194.845 27.645 195.415 ;
  END
 END i122
 PIN i123
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 199.025 27.645 199.595 ;
  END
 END i123
 PIN i124
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 203.015 27.645 203.585 ;
  END
 END i124
 PIN i125
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 207.195 27.645 207.765 ;
  END
 END i125
 PIN i126
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 19.475 27.645 20.045 ;
  END
 END i126
 PIN i127
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 211.185 27.645 211.755 ;
  END
 END i127
 PIN i128
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 215.365 27.645 215.935 ;
  END
 END i128
 PIN i129
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 237.595 27.645 238.165 ;
  END
 END i129
 PIN i130
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 241.775 27.645 242.345 ;
  END
 END i130
 PIN i131
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 245.765 27.645 246.335 ;
  END
 END i131
 PIN i132
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 249.945 27.645 250.515 ;
  END
 END i132
 PIN i133
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 253.935 27.645 254.505 ;
  END
 END i133
 PIN i134
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 258.115 27.645 258.685 ;
  END
 END i134
 PIN i135
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 262.105 27.645 262.675 ;
  END
 END i135
 PIN i136
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 266.285 27.645 266.855 ;
  END
 END i136
 PIN i137
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 23.655 27.645 24.225 ;
  END
 END i137
 PIN i138
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 270.275 27.645 270.845 ;
  END
 END i138
 PIN i139
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 274.455 27.645 275.025 ;
  END
 END i139
 PIN i140
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 278.445 27.645 279.015 ;
  END
 END i140
 PIN i141
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 282.625 27.645 283.195 ;
  END
 END i141
 PIN i142
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 286.615 27.645 287.185 ;
  END
 END i142
 PIN i143
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 27.645 27.645 28.215 ;
  END
 END i143
 PIN i144
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 31.825 27.645 32.395 ;
  END
 END i144
 PIN i145
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 35.815 27.645 36.385 ;
  END
 END i145
 PIN i146
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 39.995 27.645 40.565 ;
  END
 END i146
 PIN i147
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 142.215 3.705 142.785 ;
  END
 END i147
 PIN i148
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 142.595 4.465 143.165 ;
  END
 END i148
 PIN i149
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 3.705 28.405 4.275 ;
  END
 END i149
 PIN i150
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 7.885 28.405 8.455 ;
  END
 END i150
 PIN i151
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 44.555 28.405 45.125 ;
  END
 END i151
 PIN i152
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 48.735 28.405 49.305 ;
  END
 END i152
 PIN i153
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 52.725 28.405 53.295 ;
  END
 END i153
 PIN i154
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 56.905 28.405 57.475 ;
  END
 END i154
 PIN i155
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 79.135 28.405 79.705 ;
  END
 END i155
 PIN i156
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 83.315 28.405 83.885 ;
  END
 END i156
 PIN i157
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 87.305 28.405 87.875 ;
  END
 END i157
 PIN i158
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 91.485 28.405 92.055 ;
  END
 END i158
 PIN i159
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 95.475 28.405 96.045 ;
  END
 END i159
 PIN i160
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 99.655 28.405 100.225 ;
  END
 END i160
 PIN i161
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 11.875 28.405 12.445 ;
  END
 END i161
 PIN i162
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 103.645 28.405 104.215 ;
  END
 END i162
 PIN i163
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 107.825 28.405 108.395 ;
  END
 END i163
 PIN i164
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 111.815 28.405 112.385 ;
  END
 END i164
 PIN i165
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 115.995 28.405 116.565 ;
  END
 END i165
 PIN i166
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 119.985 28.405 120.555 ;
  END
 END i166
 PIN i167
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 124.165 28.405 124.735 ;
  END
 END i167
 PIN i168
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 128.155 28.405 128.725 ;
  END
 END i168
 PIN i169
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 132.335 28.405 132.905 ;
  END
 END i169
 PIN i170
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 161.595 28.405 162.165 ;
  END
 END i170
 PIN i171
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 165.775 28.405 166.345 ;
  END
 END i171
 PIN i172
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 16.055 28.405 16.625 ;
  END
 END i172
 PIN i173
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 169.765 28.405 170.335 ;
  END
 END i173
 PIN i174
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 173.945 28.405 174.515 ;
  END
 END i174
 PIN i175
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 177.935 28.405 178.505 ;
  END
 END i175
 PIN i176
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 182.115 28.405 182.685 ;
  END
 END i176
 PIN i177
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 186.105 28.405 186.675 ;
  END
 END i177
 PIN i178
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 190.285 28.405 190.855 ;
  END
 END i178
 PIN i179
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 194.275 28.405 194.845 ;
  END
 END i179
 PIN i180
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 198.455 28.405 199.025 ;
  END
 END i180
 PIN i181
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 202.445 28.405 203.015 ;
  END
 END i181
 PIN i182
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 206.625 28.405 207.195 ;
  END
 END i182
 PIN i183
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 20.045 28.405 20.615 ;
  END
 END i183
 PIN i184
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 210.615 28.405 211.185 ;
  END
 END i184
 PIN i185
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 214.795 28.405 215.365 ;
  END
 END i185
 PIN i186
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 237.025 28.405 237.595 ;
  END
 END i186
 PIN i187
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 241.205 28.405 241.775 ;
  END
 END i187
 PIN i188
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 245.195 28.405 245.765 ;
  END
 END i188
 PIN i189
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 249.375 28.405 249.945 ;
  END
 END i189
 PIN i190
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 253.365 28.405 253.935 ;
  END
 END i190
 PIN i191
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 257.545 28.405 258.115 ;
  END
 END i191
 PIN i192
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 261.535 28.405 262.105 ;
  END
 END i192
 PIN i193
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 265.715 28.405 266.285 ;
  END
 END i193
 PIN i194
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 24.225 28.405 24.795 ;
  END
 END i194
 PIN i195
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 269.705 28.405 270.275 ;
  END
 END i195
 PIN i196
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 273.885 28.405 274.455 ;
  END
 END i196
 PIN i197
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 277.875 28.405 278.445 ;
  END
 END i197
 PIN i198
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 282.055 28.405 282.625 ;
  END
 END i198
 PIN i199
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 286.045 28.405 286.615 ;
  END
 END i199
 PIN i200
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 28.215 28.405 28.785 ;
  END
 END i200
 PIN i201
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 32.395 28.405 32.965 ;
  END
 END i201
 PIN i202
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 36.385 28.405 36.955 ;
  END
 END i202
 PIN i203
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 40.565 28.405 41.135 ;
  END
 END i203
 PIN i204
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 4.275 134.615 4.845 135.185 ;
  END
 END i204
 PIN i205
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 5.415 134.615 5.985 135.185 ;
  END
 END i205
 PIN i206
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 6.935 134.615 7.505 135.185 ;
  END
 END i206
 PIN i207
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 8.835 134.615 9.405 135.185 ;
  END
 END i207
 PIN i208
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.975 134.615 10.545 135.185 ;
  END
 END i208
 PIN i209
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 4.275 147.915 4.845 148.485 ;
  END
 END i209
 PIN i210
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 5.415 147.915 5.985 148.485 ;
  END
 END i210
 PIN i211
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 6.935 147.915 7.505 148.485 ;
  END
 END i211
 PIN i212
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 8.835 147.915 9.405 148.485 ;
  END
 END i212
 PIN i213
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.975 147.915 10.545 148.485 ;
  END
 END i213
 OBS
  LAYER metal1 ;
   RECT 23.18 0.0 202.54 1.71 ;
   RECT 23.18 1.71 202.54 3.42 ;
   RECT 23.18 3.42 202.54 5.13 ;
   RECT 23.18 5.13 202.54 6.84 ;
   RECT 23.18 6.84 202.54 8.55 ;
   RECT 23.18 8.55 202.54 10.26 ;
   RECT 23.18 10.26 202.54 11.97 ;
   RECT 23.18 11.97 202.54 13.68 ;
   RECT 23.18 13.68 202.54 15.39 ;
   RECT 23.18 15.39 202.54 17.1 ;
   RECT 23.18 17.1 202.54 18.81 ;
   RECT 23.18 18.81 202.54 20.52 ;
   RECT 23.18 20.52 202.54 22.23 ;
   RECT 23.18 22.23 202.54 23.94 ;
   RECT 23.18 23.94 202.54 25.65 ;
   RECT 23.18 25.65 202.54 27.36 ;
   RECT 23.18 27.36 202.54 29.07 ;
   RECT 23.18 29.07 202.54 30.78 ;
   RECT 23.18 30.78 202.54 32.49 ;
   RECT 23.18 32.49 202.54 34.2 ;
   RECT 23.18 34.2 202.54 35.91 ;
   RECT 23.18 35.91 202.54 37.62 ;
   RECT 23.18 37.62 202.54 39.33 ;
   RECT 23.18 39.33 202.54 41.04 ;
   RECT 23.18 41.04 202.54 42.75 ;
   RECT 23.18 42.75 202.54 44.46 ;
   RECT 23.18 44.46 202.54 46.17 ;
   RECT 23.18 46.17 202.54 47.88 ;
   RECT 23.18 47.88 202.54 49.59 ;
   RECT 23.18 49.59 202.54 51.3 ;
   RECT 23.18 51.3 202.54 53.01 ;
   RECT 23.18 53.01 202.54 54.72 ;
   RECT 23.18 54.72 202.54 56.43 ;
   RECT 23.18 56.43 202.54 58.14 ;
   RECT 23.18 58.14 202.54 59.85 ;
   RECT 23.18 59.85 202.54 61.56 ;
   RECT 23.18 61.56 202.54 63.27 ;
   RECT 23.18 63.27 202.54 64.98 ;
   RECT 23.18 64.98 202.54 66.69 ;
   RECT 23.18 66.69 202.54 68.4 ;
   RECT 23.18 68.4 202.54 70.11 ;
   RECT 23.18 70.11 202.54 71.82 ;
   RECT 23.18 71.82 202.54 73.53 ;
   RECT 23.18 73.53 202.54 75.24 ;
   RECT 23.18 75.24 202.54 76.95 ;
   RECT 23.18 76.95 202.54 78.66 ;
   RECT 23.18 78.66 202.54 80.37 ;
   RECT 23.18 80.37 202.54 82.08 ;
   RECT 23.18 82.08 202.54 83.79 ;
   RECT 23.18 83.79 202.54 85.5 ;
   RECT 23.18 85.5 202.54 87.21 ;
   RECT 23.18 87.21 202.54 88.92 ;
   RECT 23.18 88.92 202.54 90.63 ;
   RECT 23.18 90.63 202.54 92.34 ;
   RECT 23.18 92.34 202.54 94.05 ;
   RECT 23.18 94.05 202.54 95.76 ;
   RECT 23.18 95.76 202.54 97.47 ;
   RECT 23.18 97.47 202.54 99.18 ;
   RECT 23.18 99.18 202.54 100.89 ;
   RECT 23.18 100.89 202.54 102.6 ;
   RECT 23.18 102.6 202.54 104.31 ;
   RECT 23.18 104.31 202.54 106.02 ;
   RECT 23.18 106.02 202.54 107.73 ;
   RECT 23.18 107.73 202.54 109.44 ;
   RECT 23.18 109.44 202.54 111.15 ;
   RECT 23.18 111.15 202.54 112.86 ;
   RECT 23.18 112.86 202.54 114.57 ;
   RECT 23.18 114.57 202.54 116.28 ;
   RECT 23.18 116.28 202.54 117.99 ;
   RECT 23.18 117.99 202.54 119.7 ;
   RECT 23.18 119.7 202.54 121.41 ;
   RECT 23.18 121.41 202.54 123.12 ;
   RECT 23.18 123.12 202.54 124.83 ;
   RECT 23.18 124.83 202.54 126.54 ;
   RECT 23.18 126.54 202.54 128.25 ;
   RECT 23.18 128.25 202.54 129.96 ;
   RECT 23.18 129.96 202.54 131.67 ;
   RECT 23.18 131.67 202.54 133.38 ;
   RECT 0.0 133.38 202.54 135.09 ;
   RECT 0.0 135.09 202.54 136.8 ;
   RECT 0.0 136.8 202.54 138.51 ;
   RECT 0.0 138.51 202.54 140.22 ;
   RECT 0.0 140.22 202.54 141.93 ;
   RECT 0.0 141.93 202.54 143.64 ;
   RECT 0.0 143.64 202.54 145.35 ;
   RECT 0.0 145.35 202.54 147.06 ;
   RECT 0.0 147.06 202.54 148.77 ;
   RECT 0.0 148.77 202.54 150.48 ;
   RECT 0.0 150.48 202.54 152.19 ;
   RECT 0.0 152.19 202.54 153.9 ;
   RECT 0.0 153.9 202.54 155.61 ;
   RECT 0.0 155.61 202.54 157.32 ;
   RECT 0.0 157.32 202.54 159.03 ;
   RECT 0.0 159.03 202.54 160.74 ;
   RECT 0.0 160.74 202.54 162.45 ;
   RECT 23.18 162.45 202.54 164.16 ;
   RECT 23.18 164.16 202.54 165.87 ;
   RECT 23.18 165.87 202.54 167.58 ;
   RECT 23.18 167.58 202.54 169.29 ;
   RECT 23.18 169.29 202.54 171.0 ;
   RECT 23.18 171.0 202.54 172.71 ;
   RECT 23.18 172.71 202.54 174.42 ;
   RECT 23.18 174.42 202.54 176.13 ;
   RECT 23.18 176.13 202.54 177.84 ;
   RECT 23.18 177.84 202.54 179.55 ;
   RECT 23.18 179.55 202.54 181.26 ;
   RECT 23.18 181.26 202.54 182.97 ;
   RECT 23.18 182.97 202.54 184.68 ;
   RECT 23.18 184.68 202.54 186.39 ;
   RECT 23.18 186.39 202.54 188.1 ;
   RECT 23.18 188.1 202.54 189.81 ;
   RECT 23.18 189.81 202.54 191.52 ;
   RECT 23.18 191.52 202.54 193.23 ;
   RECT 23.18 193.23 202.54 194.94 ;
   RECT 23.18 194.94 202.54 196.65 ;
   RECT 23.18 196.65 202.54 198.36 ;
   RECT 23.18 198.36 202.54 200.07 ;
   RECT 23.18 200.07 202.54 201.78 ;
   RECT 23.18 201.78 202.54 203.49 ;
   RECT 23.18 203.49 202.54 205.2 ;
   RECT 23.18 205.2 202.54 206.91 ;
   RECT 23.18 206.91 202.54 208.62 ;
   RECT 23.18 208.62 202.54 210.33 ;
   RECT 23.18 210.33 202.54 212.04 ;
   RECT 23.18 212.04 202.54 213.75 ;
   RECT 23.18 213.75 202.54 215.46 ;
   RECT 23.18 215.46 202.54 217.17 ;
   RECT 23.18 217.17 202.54 218.88 ;
   RECT 23.18 218.88 202.54 220.59 ;
   RECT 23.18 220.59 202.54 222.3 ;
   RECT 23.18 222.3 202.54 224.01 ;
   RECT 23.18 224.01 202.54 225.72 ;
   RECT 23.18 225.72 202.54 227.43 ;
   RECT 23.18 227.43 202.54 229.14 ;
   RECT 23.18 229.14 202.54 230.85 ;
   RECT 23.18 230.85 202.54 232.56 ;
   RECT 23.18 232.56 202.54 234.27 ;
   RECT 23.18 234.27 202.54 235.98 ;
   RECT 23.18 235.98 202.54 237.69 ;
   RECT 23.18 237.69 202.54 239.4 ;
   RECT 23.18 239.4 202.54 241.11 ;
   RECT 23.18 241.11 202.54 242.82 ;
   RECT 23.18 242.82 202.54 244.53 ;
   RECT 23.18 244.53 202.54 246.24 ;
   RECT 23.18 246.24 202.54 247.95 ;
   RECT 23.18 247.95 202.54 249.66 ;
   RECT 23.18 249.66 202.54 251.37 ;
   RECT 23.18 251.37 202.54 253.08 ;
   RECT 23.18 253.08 202.54 254.79 ;
   RECT 23.18 254.79 202.54 256.5 ;
   RECT 23.18 256.5 202.54 258.21 ;
   RECT 23.18 258.21 202.54 259.92 ;
   RECT 23.18 259.92 202.54 261.63 ;
   RECT 23.18 261.63 202.54 263.34 ;
   RECT 23.18 263.34 202.54 265.05 ;
   RECT 23.18 265.05 202.54 266.76 ;
   RECT 23.18 266.76 202.54 268.47 ;
   RECT 23.18 268.47 202.54 270.18 ;
   RECT 23.18 270.18 202.54 271.89 ;
   RECT 23.18 271.89 202.54 273.6 ;
   RECT 23.18 273.6 202.54 275.31 ;
   RECT 23.18 275.31 202.54 277.02 ;
   RECT 23.18 277.02 202.54 278.73 ;
   RECT 23.18 278.73 202.54 280.44 ;
   RECT 23.18 280.44 202.54 282.15 ;
   RECT 23.18 282.15 202.54 283.86 ;
   RECT 23.18 283.86 202.54 285.57 ;
   RECT 23.18 285.57 202.54 287.28 ;
   RECT 23.18 287.28 202.54 288.99 ;
   RECT 23.18 288.99 202.54 290.7 ;
   RECT 23.18 290.7 202.54 292.41 ;
  LAYER via1 ;
   RECT 23.18 0.0 202.54 1.71 ;
   RECT 23.18 1.71 202.54 3.42 ;
   RECT 23.18 3.42 202.54 5.13 ;
   RECT 23.18 5.13 202.54 6.84 ;
   RECT 23.18 6.84 202.54 8.55 ;
   RECT 23.18 8.55 202.54 10.26 ;
   RECT 23.18 10.26 202.54 11.97 ;
   RECT 23.18 11.97 202.54 13.68 ;
   RECT 23.18 13.68 202.54 15.39 ;
   RECT 23.18 15.39 202.54 17.1 ;
   RECT 23.18 17.1 202.54 18.81 ;
   RECT 23.18 18.81 202.54 20.52 ;
   RECT 23.18 20.52 202.54 22.23 ;
   RECT 23.18 22.23 202.54 23.94 ;
   RECT 23.18 23.94 202.54 25.65 ;
   RECT 23.18 25.65 202.54 27.36 ;
   RECT 23.18 27.36 202.54 29.07 ;
   RECT 23.18 29.07 202.54 30.78 ;
   RECT 23.18 30.78 202.54 32.49 ;
   RECT 23.18 32.49 202.54 34.2 ;
   RECT 23.18 34.2 202.54 35.91 ;
   RECT 23.18 35.91 202.54 37.62 ;
   RECT 23.18 37.62 202.54 39.33 ;
   RECT 23.18 39.33 202.54 41.04 ;
   RECT 23.18 41.04 202.54 42.75 ;
   RECT 23.18 42.75 202.54 44.46 ;
   RECT 23.18 44.46 202.54 46.17 ;
   RECT 23.18 46.17 202.54 47.88 ;
   RECT 23.18 47.88 202.54 49.59 ;
   RECT 23.18 49.59 202.54 51.3 ;
   RECT 23.18 51.3 202.54 53.01 ;
   RECT 23.18 53.01 202.54 54.72 ;
   RECT 23.18 54.72 202.54 56.43 ;
   RECT 23.18 56.43 202.54 58.14 ;
   RECT 23.18 58.14 202.54 59.85 ;
   RECT 23.18 59.85 202.54 61.56 ;
   RECT 23.18 61.56 202.54 63.27 ;
   RECT 23.18 63.27 202.54 64.98 ;
   RECT 23.18 64.98 202.54 66.69 ;
   RECT 23.18 66.69 202.54 68.4 ;
   RECT 23.18 68.4 202.54 70.11 ;
   RECT 23.18 70.11 202.54 71.82 ;
   RECT 23.18 71.82 202.54 73.53 ;
   RECT 23.18 73.53 202.54 75.24 ;
   RECT 23.18 75.24 202.54 76.95 ;
   RECT 23.18 76.95 202.54 78.66 ;
   RECT 23.18 78.66 202.54 80.37 ;
   RECT 23.18 80.37 202.54 82.08 ;
   RECT 23.18 82.08 202.54 83.79 ;
   RECT 23.18 83.79 202.54 85.5 ;
   RECT 23.18 85.5 202.54 87.21 ;
   RECT 23.18 87.21 202.54 88.92 ;
   RECT 23.18 88.92 202.54 90.63 ;
   RECT 23.18 90.63 202.54 92.34 ;
   RECT 23.18 92.34 202.54 94.05 ;
   RECT 23.18 94.05 202.54 95.76 ;
   RECT 23.18 95.76 202.54 97.47 ;
   RECT 23.18 97.47 202.54 99.18 ;
   RECT 23.18 99.18 202.54 100.89 ;
   RECT 23.18 100.89 202.54 102.6 ;
   RECT 23.18 102.6 202.54 104.31 ;
   RECT 23.18 104.31 202.54 106.02 ;
   RECT 23.18 106.02 202.54 107.73 ;
   RECT 23.18 107.73 202.54 109.44 ;
   RECT 23.18 109.44 202.54 111.15 ;
   RECT 23.18 111.15 202.54 112.86 ;
   RECT 23.18 112.86 202.54 114.57 ;
   RECT 23.18 114.57 202.54 116.28 ;
   RECT 23.18 116.28 202.54 117.99 ;
   RECT 23.18 117.99 202.54 119.7 ;
   RECT 23.18 119.7 202.54 121.41 ;
   RECT 23.18 121.41 202.54 123.12 ;
   RECT 23.18 123.12 202.54 124.83 ;
   RECT 23.18 124.83 202.54 126.54 ;
   RECT 23.18 126.54 202.54 128.25 ;
   RECT 23.18 128.25 202.54 129.96 ;
   RECT 23.18 129.96 202.54 131.67 ;
   RECT 23.18 131.67 202.54 133.38 ;
   RECT 0.0 133.38 202.54 135.09 ;
   RECT 0.0 135.09 202.54 136.8 ;
   RECT 0.0 136.8 202.54 138.51 ;
   RECT 0.0 138.51 202.54 140.22 ;
   RECT 0.0 140.22 202.54 141.93 ;
   RECT 0.0 141.93 202.54 143.64 ;
   RECT 0.0 143.64 202.54 145.35 ;
   RECT 0.0 145.35 202.54 147.06 ;
   RECT 0.0 147.06 202.54 148.77 ;
   RECT 0.0 148.77 202.54 150.48 ;
   RECT 0.0 150.48 202.54 152.19 ;
   RECT 0.0 152.19 202.54 153.9 ;
   RECT 0.0 153.9 202.54 155.61 ;
   RECT 0.0 155.61 202.54 157.32 ;
   RECT 0.0 157.32 202.54 159.03 ;
   RECT 0.0 159.03 202.54 160.74 ;
   RECT 0.0 160.74 202.54 162.45 ;
   RECT 23.18 162.45 202.54 164.16 ;
   RECT 23.18 164.16 202.54 165.87 ;
   RECT 23.18 165.87 202.54 167.58 ;
   RECT 23.18 167.58 202.54 169.29 ;
   RECT 23.18 169.29 202.54 171.0 ;
   RECT 23.18 171.0 202.54 172.71 ;
   RECT 23.18 172.71 202.54 174.42 ;
   RECT 23.18 174.42 202.54 176.13 ;
   RECT 23.18 176.13 202.54 177.84 ;
   RECT 23.18 177.84 202.54 179.55 ;
   RECT 23.18 179.55 202.54 181.26 ;
   RECT 23.18 181.26 202.54 182.97 ;
   RECT 23.18 182.97 202.54 184.68 ;
   RECT 23.18 184.68 202.54 186.39 ;
   RECT 23.18 186.39 202.54 188.1 ;
   RECT 23.18 188.1 202.54 189.81 ;
   RECT 23.18 189.81 202.54 191.52 ;
   RECT 23.18 191.52 202.54 193.23 ;
   RECT 23.18 193.23 202.54 194.94 ;
   RECT 23.18 194.94 202.54 196.65 ;
   RECT 23.18 196.65 202.54 198.36 ;
   RECT 23.18 198.36 202.54 200.07 ;
   RECT 23.18 200.07 202.54 201.78 ;
   RECT 23.18 201.78 202.54 203.49 ;
   RECT 23.18 203.49 202.54 205.2 ;
   RECT 23.18 205.2 202.54 206.91 ;
   RECT 23.18 206.91 202.54 208.62 ;
   RECT 23.18 208.62 202.54 210.33 ;
   RECT 23.18 210.33 202.54 212.04 ;
   RECT 23.18 212.04 202.54 213.75 ;
   RECT 23.18 213.75 202.54 215.46 ;
   RECT 23.18 215.46 202.54 217.17 ;
   RECT 23.18 217.17 202.54 218.88 ;
   RECT 23.18 218.88 202.54 220.59 ;
   RECT 23.18 220.59 202.54 222.3 ;
   RECT 23.18 222.3 202.54 224.01 ;
   RECT 23.18 224.01 202.54 225.72 ;
   RECT 23.18 225.72 202.54 227.43 ;
   RECT 23.18 227.43 202.54 229.14 ;
   RECT 23.18 229.14 202.54 230.85 ;
   RECT 23.18 230.85 202.54 232.56 ;
   RECT 23.18 232.56 202.54 234.27 ;
   RECT 23.18 234.27 202.54 235.98 ;
   RECT 23.18 235.98 202.54 237.69 ;
   RECT 23.18 237.69 202.54 239.4 ;
   RECT 23.18 239.4 202.54 241.11 ;
   RECT 23.18 241.11 202.54 242.82 ;
   RECT 23.18 242.82 202.54 244.53 ;
   RECT 23.18 244.53 202.54 246.24 ;
   RECT 23.18 246.24 202.54 247.95 ;
   RECT 23.18 247.95 202.54 249.66 ;
   RECT 23.18 249.66 202.54 251.37 ;
   RECT 23.18 251.37 202.54 253.08 ;
   RECT 23.18 253.08 202.54 254.79 ;
   RECT 23.18 254.79 202.54 256.5 ;
   RECT 23.18 256.5 202.54 258.21 ;
   RECT 23.18 258.21 202.54 259.92 ;
   RECT 23.18 259.92 202.54 261.63 ;
   RECT 23.18 261.63 202.54 263.34 ;
   RECT 23.18 263.34 202.54 265.05 ;
   RECT 23.18 265.05 202.54 266.76 ;
   RECT 23.18 266.76 202.54 268.47 ;
   RECT 23.18 268.47 202.54 270.18 ;
   RECT 23.18 270.18 202.54 271.89 ;
   RECT 23.18 271.89 202.54 273.6 ;
   RECT 23.18 273.6 202.54 275.31 ;
   RECT 23.18 275.31 202.54 277.02 ;
   RECT 23.18 277.02 202.54 278.73 ;
   RECT 23.18 278.73 202.54 280.44 ;
   RECT 23.18 280.44 202.54 282.15 ;
   RECT 23.18 282.15 202.54 283.86 ;
   RECT 23.18 283.86 202.54 285.57 ;
   RECT 23.18 285.57 202.54 287.28 ;
   RECT 23.18 287.28 202.54 288.99 ;
   RECT 23.18 288.99 202.54 290.7 ;
   RECT 23.18 290.7 202.54 292.41 ;
  LAYER metal2 ;
   RECT 23.18 0.0 202.54 1.71 ;
   RECT 23.18 1.71 202.54 3.42 ;
   RECT 23.18 3.42 202.54 5.13 ;
   RECT 23.18 5.13 202.54 6.84 ;
   RECT 23.18 6.84 202.54 8.55 ;
   RECT 23.18 8.55 202.54 10.26 ;
   RECT 23.18 10.26 202.54 11.97 ;
   RECT 23.18 11.97 202.54 13.68 ;
   RECT 23.18 13.68 202.54 15.39 ;
   RECT 23.18 15.39 202.54 17.1 ;
   RECT 23.18 17.1 202.54 18.81 ;
   RECT 23.18 18.81 202.54 20.52 ;
   RECT 23.18 20.52 202.54 22.23 ;
   RECT 23.18 22.23 202.54 23.94 ;
   RECT 23.18 23.94 202.54 25.65 ;
   RECT 23.18 25.65 202.54 27.36 ;
   RECT 23.18 27.36 202.54 29.07 ;
   RECT 23.18 29.07 202.54 30.78 ;
   RECT 23.18 30.78 202.54 32.49 ;
   RECT 23.18 32.49 202.54 34.2 ;
   RECT 23.18 34.2 202.54 35.91 ;
   RECT 23.18 35.91 202.54 37.62 ;
   RECT 23.18 37.62 202.54 39.33 ;
   RECT 23.18 39.33 202.54 41.04 ;
   RECT 23.18 41.04 202.54 42.75 ;
   RECT 23.18 42.75 202.54 44.46 ;
   RECT 23.18 44.46 202.54 46.17 ;
   RECT 23.18 46.17 202.54 47.88 ;
   RECT 23.18 47.88 202.54 49.59 ;
   RECT 23.18 49.59 202.54 51.3 ;
   RECT 23.18 51.3 202.54 53.01 ;
   RECT 23.18 53.01 202.54 54.72 ;
   RECT 23.18 54.72 202.54 56.43 ;
   RECT 23.18 56.43 202.54 58.14 ;
   RECT 23.18 58.14 202.54 59.85 ;
   RECT 23.18 59.85 202.54 61.56 ;
   RECT 23.18 61.56 202.54 63.27 ;
   RECT 23.18 63.27 202.54 64.98 ;
   RECT 23.18 64.98 202.54 66.69 ;
   RECT 23.18 66.69 202.54 68.4 ;
   RECT 23.18 68.4 202.54 70.11 ;
   RECT 23.18 70.11 202.54 71.82 ;
   RECT 23.18 71.82 202.54 73.53 ;
   RECT 23.18 73.53 202.54 75.24 ;
   RECT 23.18 75.24 202.54 76.95 ;
   RECT 23.18 76.95 202.54 78.66 ;
   RECT 23.18 78.66 202.54 80.37 ;
   RECT 23.18 80.37 202.54 82.08 ;
   RECT 23.18 82.08 202.54 83.79 ;
   RECT 23.18 83.79 202.54 85.5 ;
   RECT 23.18 85.5 202.54 87.21 ;
   RECT 23.18 87.21 202.54 88.92 ;
   RECT 23.18 88.92 202.54 90.63 ;
   RECT 23.18 90.63 202.54 92.34 ;
   RECT 23.18 92.34 202.54 94.05 ;
   RECT 23.18 94.05 202.54 95.76 ;
   RECT 23.18 95.76 202.54 97.47 ;
   RECT 23.18 97.47 202.54 99.18 ;
   RECT 23.18 99.18 202.54 100.89 ;
   RECT 23.18 100.89 202.54 102.6 ;
   RECT 23.18 102.6 202.54 104.31 ;
   RECT 23.18 104.31 202.54 106.02 ;
   RECT 23.18 106.02 202.54 107.73 ;
   RECT 23.18 107.73 202.54 109.44 ;
   RECT 23.18 109.44 202.54 111.15 ;
   RECT 23.18 111.15 202.54 112.86 ;
   RECT 23.18 112.86 202.54 114.57 ;
   RECT 23.18 114.57 202.54 116.28 ;
   RECT 23.18 116.28 202.54 117.99 ;
   RECT 23.18 117.99 202.54 119.7 ;
   RECT 23.18 119.7 202.54 121.41 ;
   RECT 23.18 121.41 202.54 123.12 ;
   RECT 23.18 123.12 202.54 124.83 ;
   RECT 23.18 124.83 202.54 126.54 ;
   RECT 23.18 126.54 202.54 128.25 ;
   RECT 23.18 128.25 202.54 129.96 ;
   RECT 23.18 129.96 202.54 131.67 ;
   RECT 23.18 131.67 202.54 133.38 ;
   RECT 0.0 133.38 202.54 135.09 ;
   RECT 0.0 135.09 202.54 136.8 ;
   RECT 0.0 136.8 202.54 138.51 ;
   RECT 0.0 138.51 202.54 140.22 ;
   RECT 0.0 140.22 202.54 141.93 ;
   RECT 0.0 141.93 202.54 143.64 ;
   RECT 0.0 143.64 202.54 145.35 ;
   RECT 0.0 145.35 202.54 147.06 ;
   RECT 0.0 147.06 202.54 148.77 ;
   RECT 0.0 148.77 202.54 150.48 ;
   RECT 0.0 150.48 202.54 152.19 ;
   RECT 0.0 152.19 202.54 153.9 ;
   RECT 0.0 153.9 202.54 155.61 ;
   RECT 0.0 155.61 202.54 157.32 ;
   RECT 0.0 157.32 202.54 159.03 ;
   RECT 0.0 159.03 202.54 160.74 ;
   RECT 0.0 160.74 202.54 162.45 ;
   RECT 23.18 162.45 202.54 164.16 ;
   RECT 23.18 164.16 202.54 165.87 ;
   RECT 23.18 165.87 202.54 167.58 ;
   RECT 23.18 167.58 202.54 169.29 ;
   RECT 23.18 169.29 202.54 171.0 ;
   RECT 23.18 171.0 202.54 172.71 ;
   RECT 23.18 172.71 202.54 174.42 ;
   RECT 23.18 174.42 202.54 176.13 ;
   RECT 23.18 176.13 202.54 177.84 ;
   RECT 23.18 177.84 202.54 179.55 ;
   RECT 23.18 179.55 202.54 181.26 ;
   RECT 23.18 181.26 202.54 182.97 ;
   RECT 23.18 182.97 202.54 184.68 ;
   RECT 23.18 184.68 202.54 186.39 ;
   RECT 23.18 186.39 202.54 188.1 ;
   RECT 23.18 188.1 202.54 189.81 ;
   RECT 23.18 189.81 202.54 191.52 ;
   RECT 23.18 191.52 202.54 193.23 ;
   RECT 23.18 193.23 202.54 194.94 ;
   RECT 23.18 194.94 202.54 196.65 ;
   RECT 23.18 196.65 202.54 198.36 ;
   RECT 23.18 198.36 202.54 200.07 ;
   RECT 23.18 200.07 202.54 201.78 ;
   RECT 23.18 201.78 202.54 203.49 ;
   RECT 23.18 203.49 202.54 205.2 ;
   RECT 23.18 205.2 202.54 206.91 ;
   RECT 23.18 206.91 202.54 208.62 ;
   RECT 23.18 208.62 202.54 210.33 ;
   RECT 23.18 210.33 202.54 212.04 ;
   RECT 23.18 212.04 202.54 213.75 ;
   RECT 23.18 213.75 202.54 215.46 ;
   RECT 23.18 215.46 202.54 217.17 ;
   RECT 23.18 217.17 202.54 218.88 ;
   RECT 23.18 218.88 202.54 220.59 ;
   RECT 23.18 220.59 202.54 222.3 ;
   RECT 23.18 222.3 202.54 224.01 ;
   RECT 23.18 224.01 202.54 225.72 ;
   RECT 23.18 225.72 202.54 227.43 ;
   RECT 23.18 227.43 202.54 229.14 ;
   RECT 23.18 229.14 202.54 230.85 ;
   RECT 23.18 230.85 202.54 232.56 ;
   RECT 23.18 232.56 202.54 234.27 ;
   RECT 23.18 234.27 202.54 235.98 ;
   RECT 23.18 235.98 202.54 237.69 ;
   RECT 23.18 237.69 202.54 239.4 ;
   RECT 23.18 239.4 202.54 241.11 ;
   RECT 23.18 241.11 202.54 242.82 ;
   RECT 23.18 242.82 202.54 244.53 ;
   RECT 23.18 244.53 202.54 246.24 ;
   RECT 23.18 246.24 202.54 247.95 ;
   RECT 23.18 247.95 202.54 249.66 ;
   RECT 23.18 249.66 202.54 251.37 ;
   RECT 23.18 251.37 202.54 253.08 ;
   RECT 23.18 253.08 202.54 254.79 ;
   RECT 23.18 254.79 202.54 256.5 ;
   RECT 23.18 256.5 202.54 258.21 ;
   RECT 23.18 258.21 202.54 259.92 ;
   RECT 23.18 259.92 202.54 261.63 ;
   RECT 23.18 261.63 202.54 263.34 ;
   RECT 23.18 263.34 202.54 265.05 ;
   RECT 23.18 265.05 202.54 266.76 ;
   RECT 23.18 266.76 202.54 268.47 ;
   RECT 23.18 268.47 202.54 270.18 ;
   RECT 23.18 270.18 202.54 271.89 ;
   RECT 23.18 271.89 202.54 273.6 ;
   RECT 23.18 273.6 202.54 275.31 ;
   RECT 23.18 275.31 202.54 277.02 ;
   RECT 23.18 277.02 202.54 278.73 ;
   RECT 23.18 278.73 202.54 280.44 ;
   RECT 23.18 280.44 202.54 282.15 ;
   RECT 23.18 282.15 202.54 283.86 ;
   RECT 23.18 283.86 202.54 285.57 ;
   RECT 23.18 285.57 202.54 287.28 ;
   RECT 23.18 287.28 202.54 288.99 ;
   RECT 23.18 288.99 202.54 290.7 ;
   RECT 23.18 290.7 202.54 292.41 ;
  LAYER via2 ;
   RECT 23.18 0.0 202.54 1.71 ;
   RECT 23.18 1.71 202.54 3.42 ;
   RECT 23.18 3.42 202.54 5.13 ;
   RECT 23.18 5.13 202.54 6.84 ;
   RECT 23.18 6.84 202.54 8.55 ;
   RECT 23.18 8.55 202.54 10.26 ;
   RECT 23.18 10.26 202.54 11.97 ;
   RECT 23.18 11.97 202.54 13.68 ;
   RECT 23.18 13.68 202.54 15.39 ;
   RECT 23.18 15.39 202.54 17.1 ;
   RECT 23.18 17.1 202.54 18.81 ;
   RECT 23.18 18.81 202.54 20.52 ;
   RECT 23.18 20.52 202.54 22.23 ;
   RECT 23.18 22.23 202.54 23.94 ;
   RECT 23.18 23.94 202.54 25.65 ;
   RECT 23.18 25.65 202.54 27.36 ;
   RECT 23.18 27.36 202.54 29.07 ;
   RECT 23.18 29.07 202.54 30.78 ;
   RECT 23.18 30.78 202.54 32.49 ;
   RECT 23.18 32.49 202.54 34.2 ;
   RECT 23.18 34.2 202.54 35.91 ;
   RECT 23.18 35.91 202.54 37.62 ;
   RECT 23.18 37.62 202.54 39.33 ;
   RECT 23.18 39.33 202.54 41.04 ;
   RECT 23.18 41.04 202.54 42.75 ;
   RECT 23.18 42.75 202.54 44.46 ;
   RECT 23.18 44.46 202.54 46.17 ;
   RECT 23.18 46.17 202.54 47.88 ;
   RECT 23.18 47.88 202.54 49.59 ;
   RECT 23.18 49.59 202.54 51.3 ;
   RECT 23.18 51.3 202.54 53.01 ;
   RECT 23.18 53.01 202.54 54.72 ;
   RECT 23.18 54.72 202.54 56.43 ;
   RECT 23.18 56.43 202.54 58.14 ;
   RECT 23.18 58.14 202.54 59.85 ;
   RECT 23.18 59.85 202.54 61.56 ;
   RECT 23.18 61.56 202.54 63.27 ;
   RECT 23.18 63.27 202.54 64.98 ;
   RECT 23.18 64.98 202.54 66.69 ;
   RECT 23.18 66.69 202.54 68.4 ;
   RECT 23.18 68.4 202.54 70.11 ;
   RECT 23.18 70.11 202.54 71.82 ;
   RECT 23.18 71.82 202.54 73.53 ;
   RECT 23.18 73.53 202.54 75.24 ;
   RECT 23.18 75.24 202.54 76.95 ;
   RECT 23.18 76.95 202.54 78.66 ;
   RECT 23.18 78.66 202.54 80.37 ;
   RECT 23.18 80.37 202.54 82.08 ;
   RECT 23.18 82.08 202.54 83.79 ;
   RECT 23.18 83.79 202.54 85.5 ;
   RECT 23.18 85.5 202.54 87.21 ;
   RECT 23.18 87.21 202.54 88.92 ;
   RECT 23.18 88.92 202.54 90.63 ;
   RECT 23.18 90.63 202.54 92.34 ;
   RECT 23.18 92.34 202.54 94.05 ;
   RECT 23.18 94.05 202.54 95.76 ;
   RECT 23.18 95.76 202.54 97.47 ;
   RECT 23.18 97.47 202.54 99.18 ;
   RECT 23.18 99.18 202.54 100.89 ;
   RECT 23.18 100.89 202.54 102.6 ;
   RECT 23.18 102.6 202.54 104.31 ;
   RECT 23.18 104.31 202.54 106.02 ;
   RECT 23.18 106.02 202.54 107.73 ;
   RECT 23.18 107.73 202.54 109.44 ;
   RECT 23.18 109.44 202.54 111.15 ;
   RECT 23.18 111.15 202.54 112.86 ;
   RECT 23.18 112.86 202.54 114.57 ;
   RECT 23.18 114.57 202.54 116.28 ;
   RECT 23.18 116.28 202.54 117.99 ;
   RECT 23.18 117.99 202.54 119.7 ;
   RECT 23.18 119.7 202.54 121.41 ;
   RECT 23.18 121.41 202.54 123.12 ;
   RECT 23.18 123.12 202.54 124.83 ;
   RECT 23.18 124.83 202.54 126.54 ;
   RECT 23.18 126.54 202.54 128.25 ;
   RECT 23.18 128.25 202.54 129.96 ;
   RECT 23.18 129.96 202.54 131.67 ;
   RECT 23.18 131.67 202.54 133.38 ;
   RECT 0.0 133.38 202.54 135.09 ;
   RECT 0.0 135.09 202.54 136.8 ;
   RECT 0.0 136.8 202.54 138.51 ;
   RECT 0.0 138.51 202.54 140.22 ;
   RECT 0.0 140.22 202.54 141.93 ;
   RECT 0.0 141.93 202.54 143.64 ;
   RECT 0.0 143.64 202.54 145.35 ;
   RECT 0.0 145.35 202.54 147.06 ;
   RECT 0.0 147.06 202.54 148.77 ;
   RECT 0.0 148.77 202.54 150.48 ;
   RECT 0.0 150.48 202.54 152.19 ;
   RECT 0.0 152.19 202.54 153.9 ;
   RECT 0.0 153.9 202.54 155.61 ;
   RECT 0.0 155.61 202.54 157.32 ;
   RECT 0.0 157.32 202.54 159.03 ;
   RECT 0.0 159.03 202.54 160.74 ;
   RECT 0.0 160.74 202.54 162.45 ;
   RECT 23.18 162.45 202.54 164.16 ;
   RECT 23.18 164.16 202.54 165.87 ;
   RECT 23.18 165.87 202.54 167.58 ;
   RECT 23.18 167.58 202.54 169.29 ;
   RECT 23.18 169.29 202.54 171.0 ;
   RECT 23.18 171.0 202.54 172.71 ;
   RECT 23.18 172.71 202.54 174.42 ;
   RECT 23.18 174.42 202.54 176.13 ;
   RECT 23.18 176.13 202.54 177.84 ;
   RECT 23.18 177.84 202.54 179.55 ;
   RECT 23.18 179.55 202.54 181.26 ;
   RECT 23.18 181.26 202.54 182.97 ;
   RECT 23.18 182.97 202.54 184.68 ;
   RECT 23.18 184.68 202.54 186.39 ;
   RECT 23.18 186.39 202.54 188.1 ;
   RECT 23.18 188.1 202.54 189.81 ;
   RECT 23.18 189.81 202.54 191.52 ;
   RECT 23.18 191.52 202.54 193.23 ;
   RECT 23.18 193.23 202.54 194.94 ;
   RECT 23.18 194.94 202.54 196.65 ;
   RECT 23.18 196.65 202.54 198.36 ;
   RECT 23.18 198.36 202.54 200.07 ;
   RECT 23.18 200.07 202.54 201.78 ;
   RECT 23.18 201.78 202.54 203.49 ;
   RECT 23.18 203.49 202.54 205.2 ;
   RECT 23.18 205.2 202.54 206.91 ;
   RECT 23.18 206.91 202.54 208.62 ;
   RECT 23.18 208.62 202.54 210.33 ;
   RECT 23.18 210.33 202.54 212.04 ;
   RECT 23.18 212.04 202.54 213.75 ;
   RECT 23.18 213.75 202.54 215.46 ;
   RECT 23.18 215.46 202.54 217.17 ;
   RECT 23.18 217.17 202.54 218.88 ;
   RECT 23.18 218.88 202.54 220.59 ;
   RECT 23.18 220.59 202.54 222.3 ;
   RECT 23.18 222.3 202.54 224.01 ;
   RECT 23.18 224.01 202.54 225.72 ;
   RECT 23.18 225.72 202.54 227.43 ;
   RECT 23.18 227.43 202.54 229.14 ;
   RECT 23.18 229.14 202.54 230.85 ;
   RECT 23.18 230.85 202.54 232.56 ;
   RECT 23.18 232.56 202.54 234.27 ;
   RECT 23.18 234.27 202.54 235.98 ;
   RECT 23.18 235.98 202.54 237.69 ;
   RECT 23.18 237.69 202.54 239.4 ;
   RECT 23.18 239.4 202.54 241.11 ;
   RECT 23.18 241.11 202.54 242.82 ;
   RECT 23.18 242.82 202.54 244.53 ;
   RECT 23.18 244.53 202.54 246.24 ;
   RECT 23.18 246.24 202.54 247.95 ;
   RECT 23.18 247.95 202.54 249.66 ;
   RECT 23.18 249.66 202.54 251.37 ;
   RECT 23.18 251.37 202.54 253.08 ;
   RECT 23.18 253.08 202.54 254.79 ;
   RECT 23.18 254.79 202.54 256.5 ;
   RECT 23.18 256.5 202.54 258.21 ;
   RECT 23.18 258.21 202.54 259.92 ;
   RECT 23.18 259.92 202.54 261.63 ;
   RECT 23.18 261.63 202.54 263.34 ;
   RECT 23.18 263.34 202.54 265.05 ;
   RECT 23.18 265.05 202.54 266.76 ;
   RECT 23.18 266.76 202.54 268.47 ;
   RECT 23.18 268.47 202.54 270.18 ;
   RECT 23.18 270.18 202.54 271.89 ;
   RECT 23.18 271.89 202.54 273.6 ;
   RECT 23.18 273.6 202.54 275.31 ;
   RECT 23.18 275.31 202.54 277.02 ;
   RECT 23.18 277.02 202.54 278.73 ;
   RECT 23.18 278.73 202.54 280.44 ;
   RECT 23.18 280.44 202.54 282.15 ;
   RECT 23.18 282.15 202.54 283.86 ;
   RECT 23.18 283.86 202.54 285.57 ;
   RECT 23.18 285.57 202.54 287.28 ;
   RECT 23.18 287.28 202.54 288.99 ;
   RECT 23.18 288.99 202.54 290.7 ;
   RECT 23.18 290.7 202.54 292.41 ;
  LAYER metal3 ;
   RECT 23.18 0.0 202.54 1.71 ;
   RECT 23.18 1.71 202.54 3.42 ;
   RECT 23.18 3.42 202.54 5.13 ;
   RECT 23.18 5.13 202.54 6.84 ;
   RECT 23.18 6.84 202.54 8.55 ;
   RECT 23.18 8.55 202.54 10.26 ;
   RECT 23.18 10.26 202.54 11.97 ;
   RECT 23.18 11.97 202.54 13.68 ;
   RECT 23.18 13.68 202.54 15.39 ;
   RECT 23.18 15.39 202.54 17.1 ;
   RECT 23.18 17.1 202.54 18.81 ;
   RECT 23.18 18.81 202.54 20.52 ;
   RECT 23.18 20.52 202.54 22.23 ;
   RECT 23.18 22.23 202.54 23.94 ;
   RECT 23.18 23.94 202.54 25.65 ;
   RECT 23.18 25.65 202.54 27.36 ;
   RECT 23.18 27.36 202.54 29.07 ;
   RECT 23.18 29.07 202.54 30.78 ;
   RECT 23.18 30.78 202.54 32.49 ;
   RECT 23.18 32.49 202.54 34.2 ;
   RECT 23.18 34.2 202.54 35.91 ;
   RECT 23.18 35.91 202.54 37.62 ;
   RECT 23.18 37.62 202.54 39.33 ;
   RECT 23.18 39.33 202.54 41.04 ;
   RECT 23.18 41.04 202.54 42.75 ;
   RECT 23.18 42.75 202.54 44.46 ;
   RECT 23.18 44.46 202.54 46.17 ;
   RECT 23.18 46.17 202.54 47.88 ;
   RECT 23.18 47.88 202.54 49.59 ;
   RECT 23.18 49.59 202.54 51.3 ;
   RECT 23.18 51.3 202.54 53.01 ;
   RECT 23.18 53.01 202.54 54.72 ;
   RECT 23.18 54.72 202.54 56.43 ;
   RECT 23.18 56.43 202.54 58.14 ;
   RECT 23.18 58.14 202.54 59.85 ;
   RECT 23.18 59.85 202.54 61.56 ;
   RECT 23.18 61.56 202.54 63.27 ;
   RECT 23.18 63.27 202.54 64.98 ;
   RECT 23.18 64.98 202.54 66.69 ;
   RECT 23.18 66.69 202.54 68.4 ;
   RECT 23.18 68.4 202.54 70.11 ;
   RECT 23.18 70.11 202.54 71.82 ;
   RECT 23.18 71.82 202.54 73.53 ;
   RECT 23.18 73.53 202.54 75.24 ;
   RECT 23.18 75.24 202.54 76.95 ;
   RECT 23.18 76.95 202.54 78.66 ;
   RECT 23.18 78.66 202.54 80.37 ;
   RECT 23.18 80.37 202.54 82.08 ;
   RECT 23.18 82.08 202.54 83.79 ;
   RECT 23.18 83.79 202.54 85.5 ;
   RECT 23.18 85.5 202.54 87.21 ;
   RECT 23.18 87.21 202.54 88.92 ;
   RECT 23.18 88.92 202.54 90.63 ;
   RECT 23.18 90.63 202.54 92.34 ;
   RECT 23.18 92.34 202.54 94.05 ;
   RECT 23.18 94.05 202.54 95.76 ;
   RECT 23.18 95.76 202.54 97.47 ;
   RECT 23.18 97.47 202.54 99.18 ;
   RECT 23.18 99.18 202.54 100.89 ;
   RECT 23.18 100.89 202.54 102.6 ;
   RECT 23.18 102.6 202.54 104.31 ;
   RECT 23.18 104.31 202.54 106.02 ;
   RECT 23.18 106.02 202.54 107.73 ;
   RECT 23.18 107.73 202.54 109.44 ;
   RECT 23.18 109.44 202.54 111.15 ;
   RECT 23.18 111.15 202.54 112.86 ;
   RECT 23.18 112.86 202.54 114.57 ;
   RECT 23.18 114.57 202.54 116.28 ;
   RECT 23.18 116.28 202.54 117.99 ;
   RECT 23.18 117.99 202.54 119.7 ;
   RECT 23.18 119.7 202.54 121.41 ;
   RECT 23.18 121.41 202.54 123.12 ;
   RECT 23.18 123.12 202.54 124.83 ;
   RECT 23.18 124.83 202.54 126.54 ;
   RECT 23.18 126.54 202.54 128.25 ;
   RECT 23.18 128.25 202.54 129.96 ;
   RECT 23.18 129.96 202.54 131.67 ;
   RECT 23.18 131.67 202.54 133.38 ;
   RECT 0.0 133.38 202.54 135.09 ;
   RECT 0.0 135.09 202.54 136.8 ;
   RECT 0.0 136.8 202.54 138.51 ;
   RECT 0.0 138.51 202.54 140.22 ;
   RECT 0.0 140.22 202.54 141.93 ;
   RECT 0.0 141.93 202.54 143.64 ;
   RECT 0.0 143.64 202.54 145.35 ;
   RECT 0.0 145.35 202.54 147.06 ;
   RECT 0.0 147.06 202.54 148.77 ;
   RECT 0.0 148.77 202.54 150.48 ;
   RECT 0.0 150.48 202.54 152.19 ;
   RECT 0.0 152.19 202.54 153.9 ;
   RECT 0.0 153.9 202.54 155.61 ;
   RECT 0.0 155.61 202.54 157.32 ;
   RECT 0.0 157.32 202.54 159.03 ;
   RECT 0.0 159.03 202.54 160.74 ;
   RECT 0.0 160.74 202.54 162.45 ;
   RECT 23.18 162.45 202.54 164.16 ;
   RECT 23.18 164.16 202.54 165.87 ;
   RECT 23.18 165.87 202.54 167.58 ;
   RECT 23.18 167.58 202.54 169.29 ;
   RECT 23.18 169.29 202.54 171.0 ;
   RECT 23.18 171.0 202.54 172.71 ;
   RECT 23.18 172.71 202.54 174.42 ;
   RECT 23.18 174.42 202.54 176.13 ;
   RECT 23.18 176.13 202.54 177.84 ;
   RECT 23.18 177.84 202.54 179.55 ;
   RECT 23.18 179.55 202.54 181.26 ;
   RECT 23.18 181.26 202.54 182.97 ;
   RECT 23.18 182.97 202.54 184.68 ;
   RECT 23.18 184.68 202.54 186.39 ;
   RECT 23.18 186.39 202.54 188.1 ;
   RECT 23.18 188.1 202.54 189.81 ;
   RECT 23.18 189.81 202.54 191.52 ;
   RECT 23.18 191.52 202.54 193.23 ;
   RECT 23.18 193.23 202.54 194.94 ;
   RECT 23.18 194.94 202.54 196.65 ;
   RECT 23.18 196.65 202.54 198.36 ;
   RECT 23.18 198.36 202.54 200.07 ;
   RECT 23.18 200.07 202.54 201.78 ;
   RECT 23.18 201.78 202.54 203.49 ;
   RECT 23.18 203.49 202.54 205.2 ;
   RECT 23.18 205.2 202.54 206.91 ;
   RECT 23.18 206.91 202.54 208.62 ;
   RECT 23.18 208.62 202.54 210.33 ;
   RECT 23.18 210.33 202.54 212.04 ;
   RECT 23.18 212.04 202.54 213.75 ;
   RECT 23.18 213.75 202.54 215.46 ;
   RECT 23.18 215.46 202.54 217.17 ;
   RECT 23.18 217.17 202.54 218.88 ;
   RECT 23.18 218.88 202.54 220.59 ;
   RECT 23.18 220.59 202.54 222.3 ;
   RECT 23.18 222.3 202.54 224.01 ;
   RECT 23.18 224.01 202.54 225.72 ;
   RECT 23.18 225.72 202.54 227.43 ;
   RECT 23.18 227.43 202.54 229.14 ;
   RECT 23.18 229.14 202.54 230.85 ;
   RECT 23.18 230.85 202.54 232.56 ;
   RECT 23.18 232.56 202.54 234.27 ;
   RECT 23.18 234.27 202.54 235.98 ;
   RECT 23.18 235.98 202.54 237.69 ;
   RECT 23.18 237.69 202.54 239.4 ;
   RECT 23.18 239.4 202.54 241.11 ;
   RECT 23.18 241.11 202.54 242.82 ;
   RECT 23.18 242.82 202.54 244.53 ;
   RECT 23.18 244.53 202.54 246.24 ;
   RECT 23.18 246.24 202.54 247.95 ;
   RECT 23.18 247.95 202.54 249.66 ;
   RECT 23.18 249.66 202.54 251.37 ;
   RECT 23.18 251.37 202.54 253.08 ;
   RECT 23.18 253.08 202.54 254.79 ;
   RECT 23.18 254.79 202.54 256.5 ;
   RECT 23.18 256.5 202.54 258.21 ;
   RECT 23.18 258.21 202.54 259.92 ;
   RECT 23.18 259.92 202.54 261.63 ;
   RECT 23.18 261.63 202.54 263.34 ;
   RECT 23.18 263.34 202.54 265.05 ;
   RECT 23.18 265.05 202.54 266.76 ;
   RECT 23.18 266.76 202.54 268.47 ;
   RECT 23.18 268.47 202.54 270.18 ;
   RECT 23.18 270.18 202.54 271.89 ;
   RECT 23.18 271.89 202.54 273.6 ;
   RECT 23.18 273.6 202.54 275.31 ;
   RECT 23.18 275.31 202.54 277.02 ;
   RECT 23.18 277.02 202.54 278.73 ;
   RECT 23.18 278.73 202.54 280.44 ;
   RECT 23.18 280.44 202.54 282.15 ;
   RECT 23.18 282.15 202.54 283.86 ;
   RECT 23.18 283.86 202.54 285.57 ;
   RECT 23.18 285.57 202.54 287.28 ;
   RECT 23.18 287.28 202.54 288.99 ;
   RECT 23.18 288.99 202.54 290.7 ;
   RECT 23.18 290.7 202.54 292.41 ;
  LAYER via3 ;
   RECT 23.18 0.0 202.54 1.71 ;
   RECT 23.18 1.71 202.54 3.42 ;
   RECT 23.18 3.42 202.54 5.13 ;
   RECT 23.18 5.13 202.54 6.84 ;
   RECT 23.18 6.84 202.54 8.55 ;
   RECT 23.18 8.55 202.54 10.26 ;
   RECT 23.18 10.26 202.54 11.97 ;
   RECT 23.18 11.97 202.54 13.68 ;
   RECT 23.18 13.68 202.54 15.39 ;
   RECT 23.18 15.39 202.54 17.1 ;
   RECT 23.18 17.1 202.54 18.81 ;
   RECT 23.18 18.81 202.54 20.52 ;
   RECT 23.18 20.52 202.54 22.23 ;
   RECT 23.18 22.23 202.54 23.94 ;
   RECT 23.18 23.94 202.54 25.65 ;
   RECT 23.18 25.65 202.54 27.36 ;
   RECT 23.18 27.36 202.54 29.07 ;
   RECT 23.18 29.07 202.54 30.78 ;
   RECT 23.18 30.78 202.54 32.49 ;
   RECT 23.18 32.49 202.54 34.2 ;
   RECT 23.18 34.2 202.54 35.91 ;
   RECT 23.18 35.91 202.54 37.62 ;
   RECT 23.18 37.62 202.54 39.33 ;
   RECT 23.18 39.33 202.54 41.04 ;
   RECT 23.18 41.04 202.54 42.75 ;
   RECT 23.18 42.75 202.54 44.46 ;
   RECT 23.18 44.46 202.54 46.17 ;
   RECT 23.18 46.17 202.54 47.88 ;
   RECT 23.18 47.88 202.54 49.59 ;
   RECT 23.18 49.59 202.54 51.3 ;
   RECT 23.18 51.3 202.54 53.01 ;
   RECT 23.18 53.01 202.54 54.72 ;
   RECT 23.18 54.72 202.54 56.43 ;
   RECT 23.18 56.43 202.54 58.14 ;
   RECT 23.18 58.14 202.54 59.85 ;
   RECT 23.18 59.85 202.54 61.56 ;
   RECT 23.18 61.56 202.54 63.27 ;
   RECT 23.18 63.27 202.54 64.98 ;
   RECT 23.18 64.98 202.54 66.69 ;
   RECT 23.18 66.69 202.54 68.4 ;
   RECT 23.18 68.4 202.54 70.11 ;
   RECT 23.18 70.11 202.54 71.82 ;
   RECT 23.18 71.82 202.54 73.53 ;
   RECT 23.18 73.53 202.54 75.24 ;
   RECT 23.18 75.24 202.54 76.95 ;
   RECT 23.18 76.95 202.54 78.66 ;
   RECT 23.18 78.66 202.54 80.37 ;
   RECT 23.18 80.37 202.54 82.08 ;
   RECT 23.18 82.08 202.54 83.79 ;
   RECT 23.18 83.79 202.54 85.5 ;
   RECT 23.18 85.5 202.54 87.21 ;
   RECT 23.18 87.21 202.54 88.92 ;
   RECT 23.18 88.92 202.54 90.63 ;
   RECT 23.18 90.63 202.54 92.34 ;
   RECT 23.18 92.34 202.54 94.05 ;
   RECT 23.18 94.05 202.54 95.76 ;
   RECT 23.18 95.76 202.54 97.47 ;
   RECT 23.18 97.47 202.54 99.18 ;
   RECT 23.18 99.18 202.54 100.89 ;
   RECT 23.18 100.89 202.54 102.6 ;
   RECT 23.18 102.6 202.54 104.31 ;
   RECT 23.18 104.31 202.54 106.02 ;
   RECT 23.18 106.02 202.54 107.73 ;
   RECT 23.18 107.73 202.54 109.44 ;
   RECT 23.18 109.44 202.54 111.15 ;
   RECT 23.18 111.15 202.54 112.86 ;
   RECT 23.18 112.86 202.54 114.57 ;
   RECT 23.18 114.57 202.54 116.28 ;
   RECT 23.18 116.28 202.54 117.99 ;
   RECT 23.18 117.99 202.54 119.7 ;
   RECT 23.18 119.7 202.54 121.41 ;
   RECT 23.18 121.41 202.54 123.12 ;
   RECT 23.18 123.12 202.54 124.83 ;
   RECT 23.18 124.83 202.54 126.54 ;
   RECT 23.18 126.54 202.54 128.25 ;
   RECT 23.18 128.25 202.54 129.96 ;
   RECT 23.18 129.96 202.54 131.67 ;
   RECT 23.18 131.67 202.54 133.38 ;
   RECT 0.0 133.38 202.54 135.09 ;
   RECT 0.0 135.09 202.54 136.8 ;
   RECT 0.0 136.8 202.54 138.51 ;
   RECT 0.0 138.51 202.54 140.22 ;
   RECT 0.0 140.22 202.54 141.93 ;
   RECT 0.0 141.93 202.54 143.64 ;
   RECT 0.0 143.64 202.54 145.35 ;
   RECT 0.0 145.35 202.54 147.06 ;
   RECT 0.0 147.06 202.54 148.77 ;
   RECT 0.0 148.77 202.54 150.48 ;
   RECT 0.0 150.48 202.54 152.19 ;
   RECT 0.0 152.19 202.54 153.9 ;
   RECT 0.0 153.9 202.54 155.61 ;
   RECT 0.0 155.61 202.54 157.32 ;
   RECT 0.0 157.32 202.54 159.03 ;
   RECT 0.0 159.03 202.54 160.74 ;
   RECT 0.0 160.74 202.54 162.45 ;
   RECT 23.18 162.45 202.54 164.16 ;
   RECT 23.18 164.16 202.54 165.87 ;
   RECT 23.18 165.87 202.54 167.58 ;
   RECT 23.18 167.58 202.54 169.29 ;
   RECT 23.18 169.29 202.54 171.0 ;
   RECT 23.18 171.0 202.54 172.71 ;
   RECT 23.18 172.71 202.54 174.42 ;
   RECT 23.18 174.42 202.54 176.13 ;
   RECT 23.18 176.13 202.54 177.84 ;
   RECT 23.18 177.84 202.54 179.55 ;
   RECT 23.18 179.55 202.54 181.26 ;
   RECT 23.18 181.26 202.54 182.97 ;
   RECT 23.18 182.97 202.54 184.68 ;
   RECT 23.18 184.68 202.54 186.39 ;
   RECT 23.18 186.39 202.54 188.1 ;
   RECT 23.18 188.1 202.54 189.81 ;
   RECT 23.18 189.81 202.54 191.52 ;
   RECT 23.18 191.52 202.54 193.23 ;
   RECT 23.18 193.23 202.54 194.94 ;
   RECT 23.18 194.94 202.54 196.65 ;
   RECT 23.18 196.65 202.54 198.36 ;
   RECT 23.18 198.36 202.54 200.07 ;
   RECT 23.18 200.07 202.54 201.78 ;
   RECT 23.18 201.78 202.54 203.49 ;
   RECT 23.18 203.49 202.54 205.2 ;
   RECT 23.18 205.2 202.54 206.91 ;
   RECT 23.18 206.91 202.54 208.62 ;
   RECT 23.18 208.62 202.54 210.33 ;
   RECT 23.18 210.33 202.54 212.04 ;
   RECT 23.18 212.04 202.54 213.75 ;
   RECT 23.18 213.75 202.54 215.46 ;
   RECT 23.18 215.46 202.54 217.17 ;
   RECT 23.18 217.17 202.54 218.88 ;
   RECT 23.18 218.88 202.54 220.59 ;
   RECT 23.18 220.59 202.54 222.3 ;
   RECT 23.18 222.3 202.54 224.01 ;
   RECT 23.18 224.01 202.54 225.72 ;
   RECT 23.18 225.72 202.54 227.43 ;
   RECT 23.18 227.43 202.54 229.14 ;
   RECT 23.18 229.14 202.54 230.85 ;
   RECT 23.18 230.85 202.54 232.56 ;
   RECT 23.18 232.56 202.54 234.27 ;
   RECT 23.18 234.27 202.54 235.98 ;
   RECT 23.18 235.98 202.54 237.69 ;
   RECT 23.18 237.69 202.54 239.4 ;
   RECT 23.18 239.4 202.54 241.11 ;
   RECT 23.18 241.11 202.54 242.82 ;
   RECT 23.18 242.82 202.54 244.53 ;
   RECT 23.18 244.53 202.54 246.24 ;
   RECT 23.18 246.24 202.54 247.95 ;
   RECT 23.18 247.95 202.54 249.66 ;
   RECT 23.18 249.66 202.54 251.37 ;
   RECT 23.18 251.37 202.54 253.08 ;
   RECT 23.18 253.08 202.54 254.79 ;
   RECT 23.18 254.79 202.54 256.5 ;
   RECT 23.18 256.5 202.54 258.21 ;
   RECT 23.18 258.21 202.54 259.92 ;
   RECT 23.18 259.92 202.54 261.63 ;
   RECT 23.18 261.63 202.54 263.34 ;
   RECT 23.18 263.34 202.54 265.05 ;
   RECT 23.18 265.05 202.54 266.76 ;
   RECT 23.18 266.76 202.54 268.47 ;
   RECT 23.18 268.47 202.54 270.18 ;
   RECT 23.18 270.18 202.54 271.89 ;
   RECT 23.18 271.89 202.54 273.6 ;
   RECT 23.18 273.6 202.54 275.31 ;
   RECT 23.18 275.31 202.54 277.02 ;
   RECT 23.18 277.02 202.54 278.73 ;
   RECT 23.18 278.73 202.54 280.44 ;
   RECT 23.18 280.44 202.54 282.15 ;
   RECT 23.18 282.15 202.54 283.86 ;
   RECT 23.18 283.86 202.54 285.57 ;
   RECT 23.18 285.57 202.54 287.28 ;
   RECT 23.18 287.28 202.54 288.99 ;
   RECT 23.18 288.99 202.54 290.7 ;
   RECT 23.18 290.7 202.54 292.41 ;
  LAYER metal4 ;
   RECT 23.18 0.0 202.54 1.71 ;
   RECT 23.18 1.71 202.54 3.42 ;
   RECT 23.18 3.42 202.54 5.13 ;
   RECT 23.18 5.13 202.54 6.84 ;
   RECT 23.18 6.84 202.54 8.55 ;
   RECT 23.18 8.55 202.54 10.26 ;
   RECT 23.18 10.26 202.54 11.97 ;
   RECT 23.18 11.97 202.54 13.68 ;
   RECT 23.18 13.68 202.54 15.39 ;
   RECT 23.18 15.39 202.54 17.1 ;
   RECT 23.18 17.1 202.54 18.81 ;
   RECT 23.18 18.81 202.54 20.52 ;
   RECT 23.18 20.52 202.54 22.23 ;
   RECT 23.18 22.23 202.54 23.94 ;
   RECT 23.18 23.94 202.54 25.65 ;
   RECT 23.18 25.65 202.54 27.36 ;
   RECT 23.18 27.36 202.54 29.07 ;
   RECT 23.18 29.07 202.54 30.78 ;
   RECT 23.18 30.78 202.54 32.49 ;
   RECT 23.18 32.49 202.54 34.2 ;
   RECT 23.18 34.2 202.54 35.91 ;
   RECT 23.18 35.91 202.54 37.62 ;
   RECT 23.18 37.62 202.54 39.33 ;
   RECT 23.18 39.33 202.54 41.04 ;
   RECT 23.18 41.04 202.54 42.75 ;
   RECT 23.18 42.75 202.54 44.46 ;
   RECT 23.18 44.46 202.54 46.17 ;
   RECT 23.18 46.17 202.54 47.88 ;
   RECT 23.18 47.88 202.54 49.59 ;
   RECT 23.18 49.59 202.54 51.3 ;
   RECT 23.18 51.3 202.54 53.01 ;
   RECT 23.18 53.01 202.54 54.72 ;
   RECT 23.18 54.72 202.54 56.43 ;
   RECT 23.18 56.43 202.54 58.14 ;
   RECT 23.18 58.14 202.54 59.85 ;
   RECT 23.18 59.85 202.54 61.56 ;
   RECT 23.18 61.56 202.54 63.27 ;
   RECT 23.18 63.27 202.54 64.98 ;
   RECT 23.18 64.98 202.54 66.69 ;
   RECT 23.18 66.69 202.54 68.4 ;
   RECT 23.18 68.4 202.54 70.11 ;
   RECT 23.18 70.11 202.54 71.82 ;
   RECT 23.18 71.82 202.54 73.53 ;
   RECT 23.18 73.53 202.54 75.24 ;
   RECT 23.18 75.24 202.54 76.95 ;
   RECT 23.18 76.95 202.54 78.66 ;
   RECT 23.18 78.66 202.54 80.37 ;
   RECT 23.18 80.37 202.54 82.08 ;
   RECT 23.18 82.08 202.54 83.79 ;
   RECT 23.18 83.79 202.54 85.5 ;
   RECT 23.18 85.5 202.54 87.21 ;
   RECT 23.18 87.21 202.54 88.92 ;
   RECT 23.18 88.92 202.54 90.63 ;
   RECT 23.18 90.63 202.54 92.34 ;
   RECT 23.18 92.34 202.54 94.05 ;
   RECT 23.18 94.05 202.54 95.76 ;
   RECT 23.18 95.76 202.54 97.47 ;
   RECT 23.18 97.47 202.54 99.18 ;
   RECT 23.18 99.18 202.54 100.89 ;
   RECT 23.18 100.89 202.54 102.6 ;
   RECT 23.18 102.6 202.54 104.31 ;
   RECT 23.18 104.31 202.54 106.02 ;
   RECT 23.18 106.02 202.54 107.73 ;
   RECT 23.18 107.73 202.54 109.44 ;
   RECT 23.18 109.44 202.54 111.15 ;
   RECT 23.18 111.15 202.54 112.86 ;
   RECT 23.18 112.86 202.54 114.57 ;
   RECT 23.18 114.57 202.54 116.28 ;
   RECT 23.18 116.28 202.54 117.99 ;
   RECT 23.18 117.99 202.54 119.7 ;
   RECT 23.18 119.7 202.54 121.41 ;
   RECT 23.18 121.41 202.54 123.12 ;
   RECT 23.18 123.12 202.54 124.83 ;
   RECT 23.18 124.83 202.54 126.54 ;
   RECT 23.18 126.54 202.54 128.25 ;
   RECT 23.18 128.25 202.54 129.96 ;
   RECT 23.18 129.96 202.54 131.67 ;
   RECT 23.18 131.67 202.54 133.38 ;
   RECT 0.0 133.38 202.54 135.09 ;
   RECT 0.0 135.09 202.54 136.8 ;
   RECT 0.0 136.8 202.54 138.51 ;
   RECT 0.0 138.51 202.54 140.22 ;
   RECT 0.0 140.22 202.54 141.93 ;
   RECT 0.0 141.93 202.54 143.64 ;
   RECT 0.0 143.64 202.54 145.35 ;
   RECT 0.0 145.35 202.54 147.06 ;
   RECT 0.0 147.06 202.54 148.77 ;
   RECT 0.0 148.77 202.54 150.48 ;
   RECT 0.0 150.48 202.54 152.19 ;
   RECT 0.0 152.19 202.54 153.9 ;
   RECT 0.0 153.9 202.54 155.61 ;
   RECT 0.0 155.61 202.54 157.32 ;
   RECT 0.0 157.32 202.54 159.03 ;
   RECT 0.0 159.03 202.54 160.74 ;
   RECT 0.0 160.74 202.54 162.45 ;
   RECT 23.18 162.45 202.54 164.16 ;
   RECT 23.18 164.16 202.54 165.87 ;
   RECT 23.18 165.87 202.54 167.58 ;
   RECT 23.18 167.58 202.54 169.29 ;
   RECT 23.18 169.29 202.54 171.0 ;
   RECT 23.18 171.0 202.54 172.71 ;
   RECT 23.18 172.71 202.54 174.42 ;
   RECT 23.18 174.42 202.54 176.13 ;
   RECT 23.18 176.13 202.54 177.84 ;
   RECT 23.18 177.84 202.54 179.55 ;
   RECT 23.18 179.55 202.54 181.26 ;
   RECT 23.18 181.26 202.54 182.97 ;
   RECT 23.18 182.97 202.54 184.68 ;
   RECT 23.18 184.68 202.54 186.39 ;
   RECT 23.18 186.39 202.54 188.1 ;
   RECT 23.18 188.1 202.54 189.81 ;
   RECT 23.18 189.81 202.54 191.52 ;
   RECT 23.18 191.52 202.54 193.23 ;
   RECT 23.18 193.23 202.54 194.94 ;
   RECT 23.18 194.94 202.54 196.65 ;
   RECT 23.18 196.65 202.54 198.36 ;
   RECT 23.18 198.36 202.54 200.07 ;
   RECT 23.18 200.07 202.54 201.78 ;
   RECT 23.18 201.78 202.54 203.49 ;
   RECT 23.18 203.49 202.54 205.2 ;
   RECT 23.18 205.2 202.54 206.91 ;
   RECT 23.18 206.91 202.54 208.62 ;
   RECT 23.18 208.62 202.54 210.33 ;
   RECT 23.18 210.33 202.54 212.04 ;
   RECT 23.18 212.04 202.54 213.75 ;
   RECT 23.18 213.75 202.54 215.46 ;
   RECT 23.18 215.46 202.54 217.17 ;
   RECT 23.18 217.17 202.54 218.88 ;
   RECT 23.18 218.88 202.54 220.59 ;
   RECT 23.18 220.59 202.54 222.3 ;
   RECT 23.18 222.3 202.54 224.01 ;
   RECT 23.18 224.01 202.54 225.72 ;
   RECT 23.18 225.72 202.54 227.43 ;
   RECT 23.18 227.43 202.54 229.14 ;
   RECT 23.18 229.14 202.54 230.85 ;
   RECT 23.18 230.85 202.54 232.56 ;
   RECT 23.18 232.56 202.54 234.27 ;
   RECT 23.18 234.27 202.54 235.98 ;
   RECT 23.18 235.98 202.54 237.69 ;
   RECT 23.18 237.69 202.54 239.4 ;
   RECT 23.18 239.4 202.54 241.11 ;
   RECT 23.18 241.11 202.54 242.82 ;
   RECT 23.18 242.82 202.54 244.53 ;
   RECT 23.18 244.53 202.54 246.24 ;
   RECT 23.18 246.24 202.54 247.95 ;
   RECT 23.18 247.95 202.54 249.66 ;
   RECT 23.18 249.66 202.54 251.37 ;
   RECT 23.18 251.37 202.54 253.08 ;
   RECT 23.18 253.08 202.54 254.79 ;
   RECT 23.18 254.79 202.54 256.5 ;
   RECT 23.18 256.5 202.54 258.21 ;
   RECT 23.18 258.21 202.54 259.92 ;
   RECT 23.18 259.92 202.54 261.63 ;
   RECT 23.18 261.63 202.54 263.34 ;
   RECT 23.18 263.34 202.54 265.05 ;
   RECT 23.18 265.05 202.54 266.76 ;
   RECT 23.18 266.76 202.54 268.47 ;
   RECT 23.18 268.47 202.54 270.18 ;
   RECT 23.18 270.18 202.54 271.89 ;
   RECT 23.18 271.89 202.54 273.6 ;
   RECT 23.18 273.6 202.54 275.31 ;
   RECT 23.18 275.31 202.54 277.02 ;
   RECT 23.18 277.02 202.54 278.73 ;
   RECT 23.18 278.73 202.54 280.44 ;
   RECT 23.18 280.44 202.54 282.15 ;
   RECT 23.18 282.15 202.54 283.86 ;
   RECT 23.18 283.86 202.54 285.57 ;
   RECT 23.18 285.57 202.54 287.28 ;
   RECT 23.18 287.28 202.54 288.99 ;
   RECT 23.18 288.99 202.54 290.7 ;
   RECT 23.18 290.7 202.54 292.41 ;
 END
END block_533x1539_269

MACRO block_671x801_111
 CLASS BLOCK ;
 FOREIGN block_671x801_111 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 254.98 BY 152.19 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 116.945 56.525 117.515 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 107.445 56.525 108.015 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 97.945 56.525 98.515 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 88.445 56.525 89.015 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 78.945 56.525 79.515 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 69.445 56.525 70.015 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 59.945 56.525 60.515 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 50.445 56.525 51.015 ;
  END
 END o7
 PIN o8
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 40.945 56.525 41.515 ;
  END
 END o8
 PIN o9
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 25.555 3.705 26.125 ;
  END
 END o9
 PIN o10
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 126.445 56.525 127.015 ;
  END
 END o10
 PIN o11
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 37.715 56.525 38.285 ;
  END
 END o11
 PIN o12
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 47.215 56.525 47.785 ;
  END
 END o12
 PIN o13
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 56.715 56.525 57.285 ;
  END
 END o13
 PIN o14
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 66.215 56.525 66.785 ;
  END
 END o14
 PIN o15
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 75.715 56.525 76.285 ;
  END
 END o15
 PIN o16
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 85.215 56.525 85.785 ;
  END
 END o16
 PIN o17
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 94.715 56.525 95.285 ;
  END
 END o17
 PIN o18
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 104.215 56.525 104.785 ;
  END
 END o18
 PIN o19
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 113.715 56.525 114.285 ;
  END
 END o19
 PIN o20
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 123.215 56.525 123.785 ;
  END
 END o20
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 16.435 3.705 17.005 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 22.325 3.705 22.895 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 16.055 4.465 16.625 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 4.655 3.705 5.225 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 6.555 3.705 7.125 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 5.605 3.705 6.175 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 18.145 3.705 18.715 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 19.095 3.705 19.665 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 13.395 3.705 13.965 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 23.275 3.705 23.845 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 101.555 56.525 102.125 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 92.055 56.525 92.625 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 82.555 56.525 83.125 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 73.055 56.525 73.625 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 63.555 56.525 64.125 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 54.055 56.525 54.625 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 111.055 56.525 111.625 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 44.555 56.525 45.125 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 35.055 56.525 35.625 ;
  END
 END i18
 PIN i19
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 120.555 56.525 121.125 ;
  END
 END i19
 PIN i20
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 0.855 3.705 1.425 ;
  END
 END i20
 PIN i21
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 26.125 4.465 26.695 ;
  END
 END i21
 PIN i22
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 127.965 56.525 128.535 ;
  END
 END i22
 PIN i23
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 56.715 128.345 57.285 128.915 ;
  END
 END i23
 PIN i24
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 130.055 56.525 130.625 ;
  END
 END i24
 PIN i25
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 128.725 56.525 129.295 ;
  END
 END i25
 PIN i26
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 56.715 129.295 57.285 129.865 ;
  END
 END i26
 PIN i27
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 30.495 3.705 31.065 ;
  END
 END i27
 PIN i28
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 28.975 3.705 29.545 ;
  END
 END i28
 PIN i29
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 2.375 3.705 2.945 ;
  END
 END i29
 PIN i30
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 1.805 4.465 2.375 ;
  END
 END i30
 PIN i31
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 29.925 4.465 30.495 ;
  END
 END i31
 PIN i32
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 28.025 3.705 28.595 ;
  END
 END i32
 PIN i33
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 2.755 4.465 3.325 ;
  END
 END i33
 PIN i34
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 4.275 4.465 4.845 ;
  END
 END i34
 PIN i35
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 3.705 3.705 4.275 ;
  END
 END i35
 PIN i36
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 4.655 29.545 5.225 30.115 ;
  END
 END i36
 PIN i37
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 13.775 4.465 14.345 ;
  END
 END i37
 PIN i38
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 18.525 4.465 19.095 ;
  END
 END i38
 PIN i39
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 17.575 4.465 18.145 ;
  END
 END i39
 PIN i40
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 23.655 4.465 24.225 ;
  END
 END i40
 PIN i41
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 24.225 3.705 24.795 ;
  END
 END i41
 PIN i42
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 5.225 4.465 5.795 ;
  END
 END i42
 PIN i43
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 6.175 4.465 6.745 ;
  END
 END i43
 PIN i44
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 7.125 4.465 7.695 ;
  END
 END i44
 PIN i45
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 10.925 3.705 11.495 ;
  END
 END i45
 PIN i46
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 22.705 4.465 23.275 ;
  END
 END i46
 PIN i47
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 26.505 3.705 27.075 ;
  END
 END i47
 PIN i48
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 4.655 1.425 5.225 1.995 ;
  END
 END i48
 PIN i49
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 33.725 56.525 34.295 ;
  END
 END i49
 PIN i50
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 43.225 56.525 43.795 ;
  END
 END i50
 PIN i51
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 52.725 56.525 53.295 ;
  END
 END i51
 PIN i52
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 62.225 56.525 62.795 ;
  END
 END i52
 PIN i53
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 71.725 56.525 72.295 ;
  END
 END i53
 PIN i54
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 81.225 56.525 81.795 ;
  END
 END i54
 PIN i55
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 90.725 56.525 91.295 ;
  END
 END i55
 PIN i56
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 100.225 56.525 100.795 ;
  END
 END i56
 PIN i57
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 109.725 56.525 110.295 ;
  END
 END i57
 PIN i58
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 119.225 56.525 119.795 ;
  END
 END i58
 PIN i59
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 38.855 56.525 39.425 ;
  END
 END i59
 PIN i60
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 48.355 56.525 48.925 ;
  END
 END i60
 PIN i61
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 57.855 56.525 58.425 ;
  END
 END i61
 PIN i62
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 67.355 56.525 67.925 ;
  END
 END i62
 PIN i63
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 76.855 56.525 77.425 ;
  END
 END i63
 PIN i64
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 86.355 56.525 86.925 ;
  END
 END i64
 PIN i65
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 95.855 56.525 96.425 ;
  END
 END i65
 PIN i66
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 105.355 56.525 105.925 ;
  END
 END i66
 PIN i67
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 114.855 56.525 115.425 ;
  END
 END i67
 PIN i68
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 124.355 56.525 124.925 ;
  END
 END i68
 PIN i69
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 56.715 130.435 57.285 131.005 ;
  END
 END i69
 PIN i70
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 39.805 56.525 40.375 ;
  END
 END i70
 PIN i71
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 49.305 56.525 49.875 ;
  END
 END i71
 PIN i72
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 58.805 56.525 59.375 ;
  END
 END i72
 PIN i73
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 68.305 56.525 68.875 ;
  END
 END i73
 PIN i74
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 77.805 56.525 78.375 ;
  END
 END i74
 PIN i75
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 87.305 56.525 87.875 ;
  END
 END i75
 PIN i76
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 96.805 56.525 97.375 ;
  END
 END i76
 PIN i77
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 106.305 56.525 106.875 ;
  END
 END i77
 PIN i78
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 115.805 56.525 116.375 ;
  END
 END i78
 PIN i79
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 125.305 56.525 125.875 ;
  END
 END i79
 PIN i80
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 56.715 34.105 57.285 34.675 ;
  END
 END i80
 PIN i81
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 56.715 43.605 57.285 44.175 ;
  END
 END i81
 PIN i82
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 56.715 53.105 57.285 53.675 ;
  END
 END i82
 PIN i83
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 56.715 62.605 57.285 63.175 ;
  END
 END i83
 PIN i84
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 56.715 72.105 57.285 72.675 ;
  END
 END i84
 PIN i85
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 56.715 81.605 57.285 82.175 ;
  END
 END i85
 PIN i86
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 56.715 91.105 57.285 91.675 ;
  END
 END i86
 PIN i87
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 56.715 100.605 57.285 101.175 ;
  END
 END i87
 PIN i88
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 56.715 110.105 57.285 110.675 ;
  END
 END i88
 PIN i89
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 56.715 119.605 57.285 120.175 ;
  END
 END i89
 OBS
  LAYER metal1 ;
   RECT 0.0 0.0 254.98 1.71 ;
   RECT 0.0 1.71 254.98 3.42 ;
   RECT 0.0 3.42 254.98 5.13 ;
   RECT 0.0 5.13 254.98 6.84 ;
   RECT 0.0 6.84 254.98 8.55 ;
   RECT 0.0 8.55 254.98 10.26 ;
   RECT 0.0 10.26 254.98 11.97 ;
   RECT 0.0 11.97 254.98 13.68 ;
   RECT 0.0 13.68 254.98 15.39 ;
   RECT 0.0 15.39 254.98 17.1 ;
   RECT 0.0 17.1 254.98 18.81 ;
   RECT 0.0 18.81 254.98 20.52 ;
   RECT 0.0 20.52 254.98 22.23 ;
   RECT 0.0 22.23 254.98 23.94 ;
   RECT 0.0 23.94 254.98 25.65 ;
   RECT 0.0 25.65 254.98 27.36 ;
   RECT 0.0 27.36 254.98 29.07 ;
   RECT 0.0 29.07 254.98 30.78 ;
   RECT 0.0 30.78 254.98 32.49 ;
   RECT 0.0 32.49 254.98 34.2 ;
   RECT 52.82 34.2 254.98 35.91 ;
   RECT 52.82 35.91 254.98 37.62 ;
   RECT 52.82 37.62 254.98 39.33 ;
   RECT 52.82 39.33 254.98 41.04 ;
   RECT 52.82 41.04 254.98 42.75 ;
   RECT 52.82 42.75 254.98 44.46 ;
   RECT 52.82 44.46 254.98 46.17 ;
   RECT 52.82 46.17 254.98 47.88 ;
   RECT 52.82 47.88 254.98 49.59 ;
   RECT 52.82 49.59 254.98 51.3 ;
   RECT 52.82 51.3 254.98 53.01 ;
   RECT 52.82 53.01 254.98 54.72 ;
   RECT 52.82 54.72 254.98 56.43 ;
   RECT 52.82 56.43 254.98 58.14 ;
   RECT 52.82 58.14 254.98 59.85 ;
   RECT 52.82 59.85 254.98 61.56 ;
   RECT 52.82 61.56 254.98 63.27 ;
   RECT 52.82 63.27 254.98 64.98 ;
   RECT 52.82 64.98 254.98 66.69 ;
   RECT 52.82 66.69 254.98 68.4 ;
   RECT 52.82 68.4 254.98 70.11 ;
   RECT 52.82 70.11 254.98 71.82 ;
   RECT 52.82 71.82 254.98 73.53 ;
   RECT 52.82 73.53 254.98 75.24 ;
   RECT 52.82 75.24 254.98 76.95 ;
   RECT 52.82 76.95 254.98 78.66 ;
   RECT 52.82 78.66 254.98 80.37 ;
   RECT 52.82 80.37 254.98 82.08 ;
   RECT 52.82 82.08 254.98 83.79 ;
   RECT 52.82 83.79 254.98 85.5 ;
   RECT 52.82 85.5 254.98 87.21 ;
   RECT 52.82 87.21 254.98 88.92 ;
   RECT 52.82 88.92 254.98 90.63 ;
   RECT 52.82 90.63 254.98 92.34 ;
   RECT 52.82 92.34 254.98 94.05 ;
   RECT 52.82 94.05 254.98 95.76 ;
   RECT 52.82 95.76 254.98 97.47 ;
   RECT 52.82 97.47 254.98 99.18 ;
   RECT 52.82 99.18 254.98 100.89 ;
   RECT 52.82 100.89 254.98 102.6 ;
   RECT 52.82 102.6 254.98 104.31 ;
   RECT 52.82 104.31 254.98 106.02 ;
   RECT 52.82 106.02 254.98 107.73 ;
   RECT 52.82 107.73 254.98 109.44 ;
   RECT 52.82 109.44 254.98 111.15 ;
   RECT 52.82 111.15 254.98 112.86 ;
   RECT 52.82 112.86 254.98 114.57 ;
   RECT 52.82 114.57 254.98 116.28 ;
   RECT 52.82 116.28 254.98 117.99 ;
   RECT 52.82 117.99 254.98 119.7 ;
   RECT 52.82 119.7 254.98 121.41 ;
   RECT 52.82 121.41 254.98 123.12 ;
   RECT 52.82 123.12 254.98 124.83 ;
   RECT 52.82 124.83 254.98 126.54 ;
   RECT 52.82 126.54 254.98 128.25 ;
   RECT 52.82 128.25 254.98 129.96 ;
   RECT 52.82 129.96 254.98 131.67 ;
   RECT 52.82 131.67 254.98 133.38 ;
   RECT 52.82 133.38 254.98 135.09 ;
   RECT 52.82 135.09 254.98 136.8 ;
   RECT 52.82 136.8 254.98 138.51 ;
   RECT 52.82 138.51 254.98 140.22 ;
   RECT 52.82 140.22 254.98 141.93 ;
   RECT 52.82 141.93 254.98 143.64 ;
   RECT 52.82 143.64 254.98 145.35 ;
   RECT 52.82 145.35 254.98 147.06 ;
   RECT 52.82 147.06 254.98 148.77 ;
   RECT 52.82 148.77 254.98 150.48 ;
   RECT 52.82 150.48 254.98 152.19 ;
  LAYER via1 ;
   RECT 0.0 0.0 254.98 1.71 ;
   RECT 0.0 1.71 254.98 3.42 ;
   RECT 0.0 3.42 254.98 5.13 ;
   RECT 0.0 5.13 254.98 6.84 ;
   RECT 0.0 6.84 254.98 8.55 ;
   RECT 0.0 8.55 254.98 10.26 ;
   RECT 0.0 10.26 254.98 11.97 ;
   RECT 0.0 11.97 254.98 13.68 ;
   RECT 0.0 13.68 254.98 15.39 ;
   RECT 0.0 15.39 254.98 17.1 ;
   RECT 0.0 17.1 254.98 18.81 ;
   RECT 0.0 18.81 254.98 20.52 ;
   RECT 0.0 20.52 254.98 22.23 ;
   RECT 0.0 22.23 254.98 23.94 ;
   RECT 0.0 23.94 254.98 25.65 ;
   RECT 0.0 25.65 254.98 27.36 ;
   RECT 0.0 27.36 254.98 29.07 ;
   RECT 0.0 29.07 254.98 30.78 ;
   RECT 0.0 30.78 254.98 32.49 ;
   RECT 0.0 32.49 254.98 34.2 ;
   RECT 52.82 34.2 254.98 35.91 ;
   RECT 52.82 35.91 254.98 37.62 ;
   RECT 52.82 37.62 254.98 39.33 ;
   RECT 52.82 39.33 254.98 41.04 ;
   RECT 52.82 41.04 254.98 42.75 ;
   RECT 52.82 42.75 254.98 44.46 ;
   RECT 52.82 44.46 254.98 46.17 ;
   RECT 52.82 46.17 254.98 47.88 ;
   RECT 52.82 47.88 254.98 49.59 ;
   RECT 52.82 49.59 254.98 51.3 ;
   RECT 52.82 51.3 254.98 53.01 ;
   RECT 52.82 53.01 254.98 54.72 ;
   RECT 52.82 54.72 254.98 56.43 ;
   RECT 52.82 56.43 254.98 58.14 ;
   RECT 52.82 58.14 254.98 59.85 ;
   RECT 52.82 59.85 254.98 61.56 ;
   RECT 52.82 61.56 254.98 63.27 ;
   RECT 52.82 63.27 254.98 64.98 ;
   RECT 52.82 64.98 254.98 66.69 ;
   RECT 52.82 66.69 254.98 68.4 ;
   RECT 52.82 68.4 254.98 70.11 ;
   RECT 52.82 70.11 254.98 71.82 ;
   RECT 52.82 71.82 254.98 73.53 ;
   RECT 52.82 73.53 254.98 75.24 ;
   RECT 52.82 75.24 254.98 76.95 ;
   RECT 52.82 76.95 254.98 78.66 ;
   RECT 52.82 78.66 254.98 80.37 ;
   RECT 52.82 80.37 254.98 82.08 ;
   RECT 52.82 82.08 254.98 83.79 ;
   RECT 52.82 83.79 254.98 85.5 ;
   RECT 52.82 85.5 254.98 87.21 ;
   RECT 52.82 87.21 254.98 88.92 ;
   RECT 52.82 88.92 254.98 90.63 ;
   RECT 52.82 90.63 254.98 92.34 ;
   RECT 52.82 92.34 254.98 94.05 ;
   RECT 52.82 94.05 254.98 95.76 ;
   RECT 52.82 95.76 254.98 97.47 ;
   RECT 52.82 97.47 254.98 99.18 ;
   RECT 52.82 99.18 254.98 100.89 ;
   RECT 52.82 100.89 254.98 102.6 ;
   RECT 52.82 102.6 254.98 104.31 ;
   RECT 52.82 104.31 254.98 106.02 ;
   RECT 52.82 106.02 254.98 107.73 ;
   RECT 52.82 107.73 254.98 109.44 ;
   RECT 52.82 109.44 254.98 111.15 ;
   RECT 52.82 111.15 254.98 112.86 ;
   RECT 52.82 112.86 254.98 114.57 ;
   RECT 52.82 114.57 254.98 116.28 ;
   RECT 52.82 116.28 254.98 117.99 ;
   RECT 52.82 117.99 254.98 119.7 ;
   RECT 52.82 119.7 254.98 121.41 ;
   RECT 52.82 121.41 254.98 123.12 ;
   RECT 52.82 123.12 254.98 124.83 ;
   RECT 52.82 124.83 254.98 126.54 ;
   RECT 52.82 126.54 254.98 128.25 ;
   RECT 52.82 128.25 254.98 129.96 ;
   RECT 52.82 129.96 254.98 131.67 ;
   RECT 52.82 131.67 254.98 133.38 ;
   RECT 52.82 133.38 254.98 135.09 ;
   RECT 52.82 135.09 254.98 136.8 ;
   RECT 52.82 136.8 254.98 138.51 ;
   RECT 52.82 138.51 254.98 140.22 ;
   RECT 52.82 140.22 254.98 141.93 ;
   RECT 52.82 141.93 254.98 143.64 ;
   RECT 52.82 143.64 254.98 145.35 ;
   RECT 52.82 145.35 254.98 147.06 ;
   RECT 52.82 147.06 254.98 148.77 ;
   RECT 52.82 148.77 254.98 150.48 ;
   RECT 52.82 150.48 254.98 152.19 ;
  LAYER metal2 ;
   RECT 0.0 0.0 254.98 1.71 ;
   RECT 0.0 1.71 254.98 3.42 ;
   RECT 0.0 3.42 254.98 5.13 ;
   RECT 0.0 5.13 254.98 6.84 ;
   RECT 0.0 6.84 254.98 8.55 ;
   RECT 0.0 8.55 254.98 10.26 ;
   RECT 0.0 10.26 254.98 11.97 ;
   RECT 0.0 11.97 254.98 13.68 ;
   RECT 0.0 13.68 254.98 15.39 ;
   RECT 0.0 15.39 254.98 17.1 ;
   RECT 0.0 17.1 254.98 18.81 ;
   RECT 0.0 18.81 254.98 20.52 ;
   RECT 0.0 20.52 254.98 22.23 ;
   RECT 0.0 22.23 254.98 23.94 ;
   RECT 0.0 23.94 254.98 25.65 ;
   RECT 0.0 25.65 254.98 27.36 ;
   RECT 0.0 27.36 254.98 29.07 ;
   RECT 0.0 29.07 254.98 30.78 ;
   RECT 0.0 30.78 254.98 32.49 ;
   RECT 0.0 32.49 254.98 34.2 ;
   RECT 52.82 34.2 254.98 35.91 ;
   RECT 52.82 35.91 254.98 37.62 ;
   RECT 52.82 37.62 254.98 39.33 ;
   RECT 52.82 39.33 254.98 41.04 ;
   RECT 52.82 41.04 254.98 42.75 ;
   RECT 52.82 42.75 254.98 44.46 ;
   RECT 52.82 44.46 254.98 46.17 ;
   RECT 52.82 46.17 254.98 47.88 ;
   RECT 52.82 47.88 254.98 49.59 ;
   RECT 52.82 49.59 254.98 51.3 ;
   RECT 52.82 51.3 254.98 53.01 ;
   RECT 52.82 53.01 254.98 54.72 ;
   RECT 52.82 54.72 254.98 56.43 ;
   RECT 52.82 56.43 254.98 58.14 ;
   RECT 52.82 58.14 254.98 59.85 ;
   RECT 52.82 59.85 254.98 61.56 ;
   RECT 52.82 61.56 254.98 63.27 ;
   RECT 52.82 63.27 254.98 64.98 ;
   RECT 52.82 64.98 254.98 66.69 ;
   RECT 52.82 66.69 254.98 68.4 ;
   RECT 52.82 68.4 254.98 70.11 ;
   RECT 52.82 70.11 254.98 71.82 ;
   RECT 52.82 71.82 254.98 73.53 ;
   RECT 52.82 73.53 254.98 75.24 ;
   RECT 52.82 75.24 254.98 76.95 ;
   RECT 52.82 76.95 254.98 78.66 ;
   RECT 52.82 78.66 254.98 80.37 ;
   RECT 52.82 80.37 254.98 82.08 ;
   RECT 52.82 82.08 254.98 83.79 ;
   RECT 52.82 83.79 254.98 85.5 ;
   RECT 52.82 85.5 254.98 87.21 ;
   RECT 52.82 87.21 254.98 88.92 ;
   RECT 52.82 88.92 254.98 90.63 ;
   RECT 52.82 90.63 254.98 92.34 ;
   RECT 52.82 92.34 254.98 94.05 ;
   RECT 52.82 94.05 254.98 95.76 ;
   RECT 52.82 95.76 254.98 97.47 ;
   RECT 52.82 97.47 254.98 99.18 ;
   RECT 52.82 99.18 254.98 100.89 ;
   RECT 52.82 100.89 254.98 102.6 ;
   RECT 52.82 102.6 254.98 104.31 ;
   RECT 52.82 104.31 254.98 106.02 ;
   RECT 52.82 106.02 254.98 107.73 ;
   RECT 52.82 107.73 254.98 109.44 ;
   RECT 52.82 109.44 254.98 111.15 ;
   RECT 52.82 111.15 254.98 112.86 ;
   RECT 52.82 112.86 254.98 114.57 ;
   RECT 52.82 114.57 254.98 116.28 ;
   RECT 52.82 116.28 254.98 117.99 ;
   RECT 52.82 117.99 254.98 119.7 ;
   RECT 52.82 119.7 254.98 121.41 ;
   RECT 52.82 121.41 254.98 123.12 ;
   RECT 52.82 123.12 254.98 124.83 ;
   RECT 52.82 124.83 254.98 126.54 ;
   RECT 52.82 126.54 254.98 128.25 ;
   RECT 52.82 128.25 254.98 129.96 ;
   RECT 52.82 129.96 254.98 131.67 ;
   RECT 52.82 131.67 254.98 133.38 ;
   RECT 52.82 133.38 254.98 135.09 ;
   RECT 52.82 135.09 254.98 136.8 ;
   RECT 52.82 136.8 254.98 138.51 ;
   RECT 52.82 138.51 254.98 140.22 ;
   RECT 52.82 140.22 254.98 141.93 ;
   RECT 52.82 141.93 254.98 143.64 ;
   RECT 52.82 143.64 254.98 145.35 ;
   RECT 52.82 145.35 254.98 147.06 ;
   RECT 52.82 147.06 254.98 148.77 ;
   RECT 52.82 148.77 254.98 150.48 ;
   RECT 52.82 150.48 254.98 152.19 ;
  LAYER via2 ;
   RECT 0.0 0.0 254.98 1.71 ;
   RECT 0.0 1.71 254.98 3.42 ;
   RECT 0.0 3.42 254.98 5.13 ;
   RECT 0.0 5.13 254.98 6.84 ;
   RECT 0.0 6.84 254.98 8.55 ;
   RECT 0.0 8.55 254.98 10.26 ;
   RECT 0.0 10.26 254.98 11.97 ;
   RECT 0.0 11.97 254.98 13.68 ;
   RECT 0.0 13.68 254.98 15.39 ;
   RECT 0.0 15.39 254.98 17.1 ;
   RECT 0.0 17.1 254.98 18.81 ;
   RECT 0.0 18.81 254.98 20.52 ;
   RECT 0.0 20.52 254.98 22.23 ;
   RECT 0.0 22.23 254.98 23.94 ;
   RECT 0.0 23.94 254.98 25.65 ;
   RECT 0.0 25.65 254.98 27.36 ;
   RECT 0.0 27.36 254.98 29.07 ;
   RECT 0.0 29.07 254.98 30.78 ;
   RECT 0.0 30.78 254.98 32.49 ;
   RECT 0.0 32.49 254.98 34.2 ;
   RECT 52.82 34.2 254.98 35.91 ;
   RECT 52.82 35.91 254.98 37.62 ;
   RECT 52.82 37.62 254.98 39.33 ;
   RECT 52.82 39.33 254.98 41.04 ;
   RECT 52.82 41.04 254.98 42.75 ;
   RECT 52.82 42.75 254.98 44.46 ;
   RECT 52.82 44.46 254.98 46.17 ;
   RECT 52.82 46.17 254.98 47.88 ;
   RECT 52.82 47.88 254.98 49.59 ;
   RECT 52.82 49.59 254.98 51.3 ;
   RECT 52.82 51.3 254.98 53.01 ;
   RECT 52.82 53.01 254.98 54.72 ;
   RECT 52.82 54.72 254.98 56.43 ;
   RECT 52.82 56.43 254.98 58.14 ;
   RECT 52.82 58.14 254.98 59.85 ;
   RECT 52.82 59.85 254.98 61.56 ;
   RECT 52.82 61.56 254.98 63.27 ;
   RECT 52.82 63.27 254.98 64.98 ;
   RECT 52.82 64.98 254.98 66.69 ;
   RECT 52.82 66.69 254.98 68.4 ;
   RECT 52.82 68.4 254.98 70.11 ;
   RECT 52.82 70.11 254.98 71.82 ;
   RECT 52.82 71.82 254.98 73.53 ;
   RECT 52.82 73.53 254.98 75.24 ;
   RECT 52.82 75.24 254.98 76.95 ;
   RECT 52.82 76.95 254.98 78.66 ;
   RECT 52.82 78.66 254.98 80.37 ;
   RECT 52.82 80.37 254.98 82.08 ;
   RECT 52.82 82.08 254.98 83.79 ;
   RECT 52.82 83.79 254.98 85.5 ;
   RECT 52.82 85.5 254.98 87.21 ;
   RECT 52.82 87.21 254.98 88.92 ;
   RECT 52.82 88.92 254.98 90.63 ;
   RECT 52.82 90.63 254.98 92.34 ;
   RECT 52.82 92.34 254.98 94.05 ;
   RECT 52.82 94.05 254.98 95.76 ;
   RECT 52.82 95.76 254.98 97.47 ;
   RECT 52.82 97.47 254.98 99.18 ;
   RECT 52.82 99.18 254.98 100.89 ;
   RECT 52.82 100.89 254.98 102.6 ;
   RECT 52.82 102.6 254.98 104.31 ;
   RECT 52.82 104.31 254.98 106.02 ;
   RECT 52.82 106.02 254.98 107.73 ;
   RECT 52.82 107.73 254.98 109.44 ;
   RECT 52.82 109.44 254.98 111.15 ;
   RECT 52.82 111.15 254.98 112.86 ;
   RECT 52.82 112.86 254.98 114.57 ;
   RECT 52.82 114.57 254.98 116.28 ;
   RECT 52.82 116.28 254.98 117.99 ;
   RECT 52.82 117.99 254.98 119.7 ;
   RECT 52.82 119.7 254.98 121.41 ;
   RECT 52.82 121.41 254.98 123.12 ;
   RECT 52.82 123.12 254.98 124.83 ;
   RECT 52.82 124.83 254.98 126.54 ;
   RECT 52.82 126.54 254.98 128.25 ;
   RECT 52.82 128.25 254.98 129.96 ;
   RECT 52.82 129.96 254.98 131.67 ;
   RECT 52.82 131.67 254.98 133.38 ;
   RECT 52.82 133.38 254.98 135.09 ;
   RECT 52.82 135.09 254.98 136.8 ;
   RECT 52.82 136.8 254.98 138.51 ;
   RECT 52.82 138.51 254.98 140.22 ;
   RECT 52.82 140.22 254.98 141.93 ;
   RECT 52.82 141.93 254.98 143.64 ;
   RECT 52.82 143.64 254.98 145.35 ;
   RECT 52.82 145.35 254.98 147.06 ;
   RECT 52.82 147.06 254.98 148.77 ;
   RECT 52.82 148.77 254.98 150.48 ;
   RECT 52.82 150.48 254.98 152.19 ;
  LAYER metal3 ;
   RECT 0.0 0.0 254.98 1.71 ;
   RECT 0.0 1.71 254.98 3.42 ;
   RECT 0.0 3.42 254.98 5.13 ;
   RECT 0.0 5.13 254.98 6.84 ;
   RECT 0.0 6.84 254.98 8.55 ;
   RECT 0.0 8.55 254.98 10.26 ;
   RECT 0.0 10.26 254.98 11.97 ;
   RECT 0.0 11.97 254.98 13.68 ;
   RECT 0.0 13.68 254.98 15.39 ;
   RECT 0.0 15.39 254.98 17.1 ;
   RECT 0.0 17.1 254.98 18.81 ;
   RECT 0.0 18.81 254.98 20.52 ;
   RECT 0.0 20.52 254.98 22.23 ;
   RECT 0.0 22.23 254.98 23.94 ;
   RECT 0.0 23.94 254.98 25.65 ;
   RECT 0.0 25.65 254.98 27.36 ;
   RECT 0.0 27.36 254.98 29.07 ;
   RECT 0.0 29.07 254.98 30.78 ;
   RECT 0.0 30.78 254.98 32.49 ;
   RECT 0.0 32.49 254.98 34.2 ;
   RECT 52.82 34.2 254.98 35.91 ;
   RECT 52.82 35.91 254.98 37.62 ;
   RECT 52.82 37.62 254.98 39.33 ;
   RECT 52.82 39.33 254.98 41.04 ;
   RECT 52.82 41.04 254.98 42.75 ;
   RECT 52.82 42.75 254.98 44.46 ;
   RECT 52.82 44.46 254.98 46.17 ;
   RECT 52.82 46.17 254.98 47.88 ;
   RECT 52.82 47.88 254.98 49.59 ;
   RECT 52.82 49.59 254.98 51.3 ;
   RECT 52.82 51.3 254.98 53.01 ;
   RECT 52.82 53.01 254.98 54.72 ;
   RECT 52.82 54.72 254.98 56.43 ;
   RECT 52.82 56.43 254.98 58.14 ;
   RECT 52.82 58.14 254.98 59.85 ;
   RECT 52.82 59.85 254.98 61.56 ;
   RECT 52.82 61.56 254.98 63.27 ;
   RECT 52.82 63.27 254.98 64.98 ;
   RECT 52.82 64.98 254.98 66.69 ;
   RECT 52.82 66.69 254.98 68.4 ;
   RECT 52.82 68.4 254.98 70.11 ;
   RECT 52.82 70.11 254.98 71.82 ;
   RECT 52.82 71.82 254.98 73.53 ;
   RECT 52.82 73.53 254.98 75.24 ;
   RECT 52.82 75.24 254.98 76.95 ;
   RECT 52.82 76.95 254.98 78.66 ;
   RECT 52.82 78.66 254.98 80.37 ;
   RECT 52.82 80.37 254.98 82.08 ;
   RECT 52.82 82.08 254.98 83.79 ;
   RECT 52.82 83.79 254.98 85.5 ;
   RECT 52.82 85.5 254.98 87.21 ;
   RECT 52.82 87.21 254.98 88.92 ;
   RECT 52.82 88.92 254.98 90.63 ;
   RECT 52.82 90.63 254.98 92.34 ;
   RECT 52.82 92.34 254.98 94.05 ;
   RECT 52.82 94.05 254.98 95.76 ;
   RECT 52.82 95.76 254.98 97.47 ;
   RECT 52.82 97.47 254.98 99.18 ;
   RECT 52.82 99.18 254.98 100.89 ;
   RECT 52.82 100.89 254.98 102.6 ;
   RECT 52.82 102.6 254.98 104.31 ;
   RECT 52.82 104.31 254.98 106.02 ;
   RECT 52.82 106.02 254.98 107.73 ;
   RECT 52.82 107.73 254.98 109.44 ;
   RECT 52.82 109.44 254.98 111.15 ;
   RECT 52.82 111.15 254.98 112.86 ;
   RECT 52.82 112.86 254.98 114.57 ;
   RECT 52.82 114.57 254.98 116.28 ;
   RECT 52.82 116.28 254.98 117.99 ;
   RECT 52.82 117.99 254.98 119.7 ;
   RECT 52.82 119.7 254.98 121.41 ;
   RECT 52.82 121.41 254.98 123.12 ;
   RECT 52.82 123.12 254.98 124.83 ;
   RECT 52.82 124.83 254.98 126.54 ;
   RECT 52.82 126.54 254.98 128.25 ;
   RECT 52.82 128.25 254.98 129.96 ;
   RECT 52.82 129.96 254.98 131.67 ;
   RECT 52.82 131.67 254.98 133.38 ;
   RECT 52.82 133.38 254.98 135.09 ;
   RECT 52.82 135.09 254.98 136.8 ;
   RECT 52.82 136.8 254.98 138.51 ;
   RECT 52.82 138.51 254.98 140.22 ;
   RECT 52.82 140.22 254.98 141.93 ;
   RECT 52.82 141.93 254.98 143.64 ;
   RECT 52.82 143.64 254.98 145.35 ;
   RECT 52.82 145.35 254.98 147.06 ;
   RECT 52.82 147.06 254.98 148.77 ;
   RECT 52.82 148.77 254.98 150.48 ;
   RECT 52.82 150.48 254.98 152.19 ;
  LAYER via3 ;
   RECT 0.0 0.0 254.98 1.71 ;
   RECT 0.0 1.71 254.98 3.42 ;
   RECT 0.0 3.42 254.98 5.13 ;
   RECT 0.0 5.13 254.98 6.84 ;
   RECT 0.0 6.84 254.98 8.55 ;
   RECT 0.0 8.55 254.98 10.26 ;
   RECT 0.0 10.26 254.98 11.97 ;
   RECT 0.0 11.97 254.98 13.68 ;
   RECT 0.0 13.68 254.98 15.39 ;
   RECT 0.0 15.39 254.98 17.1 ;
   RECT 0.0 17.1 254.98 18.81 ;
   RECT 0.0 18.81 254.98 20.52 ;
   RECT 0.0 20.52 254.98 22.23 ;
   RECT 0.0 22.23 254.98 23.94 ;
   RECT 0.0 23.94 254.98 25.65 ;
   RECT 0.0 25.65 254.98 27.36 ;
   RECT 0.0 27.36 254.98 29.07 ;
   RECT 0.0 29.07 254.98 30.78 ;
   RECT 0.0 30.78 254.98 32.49 ;
   RECT 0.0 32.49 254.98 34.2 ;
   RECT 52.82 34.2 254.98 35.91 ;
   RECT 52.82 35.91 254.98 37.62 ;
   RECT 52.82 37.62 254.98 39.33 ;
   RECT 52.82 39.33 254.98 41.04 ;
   RECT 52.82 41.04 254.98 42.75 ;
   RECT 52.82 42.75 254.98 44.46 ;
   RECT 52.82 44.46 254.98 46.17 ;
   RECT 52.82 46.17 254.98 47.88 ;
   RECT 52.82 47.88 254.98 49.59 ;
   RECT 52.82 49.59 254.98 51.3 ;
   RECT 52.82 51.3 254.98 53.01 ;
   RECT 52.82 53.01 254.98 54.72 ;
   RECT 52.82 54.72 254.98 56.43 ;
   RECT 52.82 56.43 254.98 58.14 ;
   RECT 52.82 58.14 254.98 59.85 ;
   RECT 52.82 59.85 254.98 61.56 ;
   RECT 52.82 61.56 254.98 63.27 ;
   RECT 52.82 63.27 254.98 64.98 ;
   RECT 52.82 64.98 254.98 66.69 ;
   RECT 52.82 66.69 254.98 68.4 ;
   RECT 52.82 68.4 254.98 70.11 ;
   RECT 52.82 70.11 254.98 71.82 ;
   RECT 52.82 71.82 254.98 73.53 ;
   RECT 52.82 73.53 254.98 75.24 ;
   RECT 52.82 75.24 254.98 76.95 ;
   RECT 52.82 76.95 254.98 78.66 ;
   RECT 52.82 78.66 254.98 80.37 ;
   RECT 52.82 80.37 254.98 82.08 ;
   RECT 52.82 82.08 254.98 83.79 ;
   RECT 52.82 83.79 254.98 85.5 ;
   RECT 52.82 85.5 254.98 87.21 ;
   RECT 52.82 87.21 254.98 88.92 ;
   RECT 52.82 88.92 254.98 90.63 ;
   RECT 52.82 90.63 254.98 92.34 ;
   RECT 52.82 92.34 254.98 94.05 ;
   RECT 52.82 94.05 254.98 95.76 ;
   RECT 52.82 95.76 254.98 97.47 ;
   RECT 52.82 97.47 254.98 99.18 ;
   RECT 52.82 99.18 254.98 100.89 ;
   RECT 52.82 100.89 254.98 102.6 ;
   RECT 52.82 102.6 254.98 104.31 ;
   RECT 52.82 104.31 254.98 106.02 ;
   RECT 52.82 106.02 254.98 107.73 ;
   RECT 52.82 107.73 254.98 109.44 ;
   RECT 52.82 109.44 254.98 111.15 ;
   RECT 52.82 111.15 254.98 112.86 ;
   RECT 52.82 112.86 254.98 114.57 ;
   RECT 52.82 114.57 254.98 116.28 ;
   RECT 52.82 116.28 254.98 117.99 ;
   RECT 52.82 117.99 254.98 119.7 ;
   RECT 52.82 119.7 254.98 121.41 ;
   RECT 52.82 121.41 254.98 123.12 ;
   RECT 52.82 123.12 254.98 124.83 ;
   RECT 52.82 124.83 254.98 126.54 ;
   RECT 52.82 126.54 254.98 128.25 ;
   RECT 52.82 128.25 254.98 129.96 ;
   RECT 52.82 129.96 254.98 131.67 ;
   RECT 52.82 131.67 254.98 133.38 ;
   RECT 52.82 133.38 254.98 135.09 ;
   RECT 52.82 135.09 254.98 136.8 ;
   RECT 52.82 136.8 254.98 138.51 ;
   RECT 52.82 138.51 254.98 140.22 ;
   RECT 52.82 140.22 254.98 141.93 ;
   RECT 52.82 141.93 254.98 143.64 ;
   RECT 52.82 143.64 254.98 145.35 ;
   RECT 52.82 145.35 254.98 147.06 ;
   RECT 52.82 147.06 254.98 148.77 ;
   RECT 52.82 148.77 254.98 150.48 ;
   RECT 52.82 150.48 254.98 152.19 ;
  LAYER metal4 ;
   RECT 0.0 0.0 254.98 1.71 ;
   RECT 0.0 1.71 254.98 3.42 ;
   RECT 0.0 3.42 254.98 5.13 ;
   RECT 0.0 5.13 254.98 6.84 ;
   RECT 0.0 6.84 254.98 8.55 ;
   RECT 0.0 8.55 254.98 10.26 ;
   RECT 0.0 10.26 254.98 11.97 ;
   RECT 0.0 11.97 254.98 13.68 ;
   RECT 0.0 13.68 254.98 15.39 ;
   RECT 0.0 15.39 254.98 17.1 ;
   RECT 0.0 17.1 254.98 18.81 ;
   RECT 0.0 18.81 254.98 20.52 ;
   RECT 0.0 20.52 254.98 22.23 ;
   RECT 0.0 22.23 254.98 23.94 ;
   RECT 0.0 23.94 254.98 25.65 ;
   RECT 0.0 25.65 254.98 27.36 ;
   RECT 0.0 27.36 254.98 29.07 ;
   RECT 0.0 29.07 254.98 30.78 ;
   RECT 0.0 30.78 254.98 32.49 ;
   RECT 0.0 32.49 254.98 34.2 ;
   RECT 52.82 34.2 254.98 35.91 ;
   RECT 52.82 35.91 254.98 37.62 ;
   RECT 52.82 37.62 254.98 39.33 ;
   RECT 52.82 39.33 254.98 41.04 ;
   RECT 52.82 41.04 254.98 42.75 ;
   RECT 52.82 42.75 254.98 44.46 ;
   RECT 52.82 44.46 254.98 46.17 ;
   RECT 52.82 46.17 254.98 47.88 ;
   RECT 52.82 47.88 254.98 49.59 ;
   RECT 52.82 49.59 254.98 51.3 ;
   RECT 52.82 51.3 254.98 53.01 ;
   RECT 52.82 53.01 254.98 54.72 ;
   RECT 52.82 54.72 254.98 56.43 ;
   RECT 52.82 56.43 254.98 58.14 ;
   RECT 52.82 58.14 254.98 59.85 ;
   RECT 52.82 59.85 254.98 61.56 ;
   RECT 52.82 61.56 254.98 63.27 ;
   RECT 52.82 63.27 254.98 64.98 ;
   RECT 52.82 64.98 254.98 66.69 ;
   RECT 52.82 66.69 254.98 68.4 ;
   RECT 52.82 68.4 254.98 70.11 ;
   RECT 52.82 70.11 254.98 71.82 ;
   RECT 52.82 71.82 254.98 73.53 ;
   RECT 52.82 73.53 254.98 75.24 ;
   RECT 52.82 75.24 254.98 76.95 ;
   RECT 52.82 76.95 254.98 78.66 ;
   RECT 52.82 78.66 254.98 80.37 ;
   RECT 52.82 80.37 254.98 82.08 ;
   RECT 52.82 82.08 254.98 83.79 ;
   RECT 52.82 83.79 254.98 85.5 ;
   RECT 52.82 85.5 254.98 87.21 ;
   RECT 52.82 87.21 254.98 88.92 ;
   RECT 52.82 88.92 254.98 90.63 ;
   RECT 52.82 90.63 254.98 92.34 ;
   RECT 52.82 92.34 254.98 94.05 ;
   RECT 52.82 94.05 254.98 95.76 ;
   RECT 52.82 95.76 254.98 97.47 ;
   RECT 52.82 97.47 254.98 99.18 ;
   RECT 52.82 99.18 254.98 100.89 ;
   RECT 52.82 100.89 254.98 102.6 ;
   RECT 52.82 102.6 254.98 104.31 ;
   RECT 52.82 104.31 254.98 106.02 ;
   RECT 52.82 106.02 254.98 107.73 ;
   RECT 52.82 107.73 254.98 109.44 ;
   RECT 52.82 109.44 254.98 111.15 ;
   RECT 52.82 111.15 254.98 112.86 ;
   RECT 52.82 112.86 254.98 114.57 ;
   RECT 52.82 114.57 254.98 116.28 ;
   RECT 52.82 116.28 254.98 117.99 ;
   RECT 52.82 117.99 254.98 119.7 ;
   RECT 52.82 119.7 254.98 121.41 ;
   RECT 52.82 121.41 254.98 123.12 ;
   RECT 52.82 123.12 254.98 124.83 ;
   RECT 52.82 124.83 254.98 126.54 ;
   RECT 52.82 126.54 254.98 128.25 ;
   RECT 52.82 128.25 254.98 129.96 ;
   RECT 52.82 129.96 254.98 131.67 ;
   RECT 52.82 131.67 254.98 133.38 ;
   RECT 52.82 133.38 254.98 135.09 ;
   RECT 52.82 135.09 254.98 136.8 ;
   RECT 52.82 136.8 254.98 138.51 ;
   RECT 52.82 138.51 254.98 140.22 ;
   RECT 52.82 140.22 254.98 141.93 ;
   RECT 52.82 141.93 254.98 143.64 ;
   RECT 52.82 143.64 254.98 145.35 ;
   RECT 52.82 145.35 254.98 147.06 ;
   RECT 52.82 147.06 254.98 148.77 ;
   RECT 52.82 148.77 254.98 150.48 ;
   RECT 52.82 150.48 254.98 152.19 ;
 END
END block_671x801_111

MACRO block_197x180_33
 CLASS BLOCK ;
 FOREIGN block_197x180_33 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 74.86 BY 34.2 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 25.175 71.725 25.745 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 16.815 71.725 17.385 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 15.295 3.325 15.865 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 16.055 3.325 16.625 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 16.815 3.325 17.385 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 17.575 3.325 18.145 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 18.335 3.325 18.905 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 12.635 3.325 13.205 ;
  END
 END o7
 PIN o8
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 18.335 71.725 18.905 ;
  END
 END o8
 PIN o9
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 9.595 3.325 10.165 ;
  END
 END o9
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 21.375 71.725 21.945 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 70.395 21.755 70.965 22.325 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 22.135 71.725 22.705 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 70.395 22.515 70.965 23.085 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 24.415 71.725 24.985 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 70.395 24.795 70.965 25.365 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 26.695 71.725 27.265 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 27.455 71.725 28.025 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 5.035 3.325 5.605 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 16.055 71.725 16.625 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 13.775 71.725 14.345 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 12.255 71.725 12.825 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 28.975 71.725 29.545 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 25.935 71.725 26.505 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 17.575 71.725 18.145 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 29.735 3.325 30.305 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 22.895 71.725 23.465 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 4.275 71.725 4.845 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 5.035 71.725 5.605 ;
  END
 END i18
 PIN i19
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 6.935 71.725 7.505 ;
  END
 END i19
 PIN i20
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 7.695 71.725 8.265 ;
  END
 END i20
 PIN i21
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 8.835 71.725 9.405 ;
  END
 END i21
 PIN i22
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 9.595 71.725 10.165 ;
  END
 END i22
 OBS
  LAYER metal1 ;
   RECT 0 0 74.86 34.2 ;
  LAYER via1 ;
   RECT 0 0 74.86 34.2 ;
  LAYER metal2 ;
   RECT 0 0 74.86 34.2 ;
  LAYER via2 ;
   RECT 0 0 74.86 34.2 ;
  LAYER metal3 ;
   RECT 0 0 74.86 34.2 ;
  LAYER via3 ;
   RECT 0 0 74.86 34.2 ;
  LAYER metal4 ;
   RECT 0 0 74.86 34.2 ;
 END
END block_197x180_33

MACRO block_1338x2160_145
 CLASS BLOCK ;
 FOREIGN block_1338x2160_145 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 508.44 BY 410.4 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 400.045 26.885 400.615 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 383.705 26.885 384.275 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 218.405 26.885 218.975 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 173.945 26.885 174.515 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 157.605 26.885 158.175 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 141.265 26.885 141.835 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 124.925 26.885 125.495 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 108.585 26.885 109.155 ;
  END
 END o7
 PIN o8
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 74.005 26.885 74.575 ;
  END
 END o8
 PIN o9
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 57.665 26.885 58.235 ;
  END
 END o9
 PIN o10
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 41.325 26.885 41.895 ;
  END
 END o10
 PIN o11
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 24.985 26.885 25.555 ;
  END
 END o11
 PIN o12
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 367.365 26.885 367.935 ;
  END
 END o12
 PIN o13
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 8.645 26.885 9.215 ;
  END
 END o13
 PIN o14
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 351.025 26.885 351.595 ;
  END
 END o14
 PIN o15
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 334.685 26.885 335.255 ;
  END
 END o15
 PIN o16
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 318.345 26.885 318.915 ;
  END
 END o16
 PIN o17
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 283.765 26.885 284.335 ;
  END
 END o17
 PIN o18
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 267.425 26.885 267.995 ;
  END
 END o18
 PIN o19
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 251.085 26.885 251.655 ;
  END
 END o19
 PIN o20
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 234.745 26.885 235.315 ;
  END
 END o20
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 207.385 3.705 207.955 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 185.725 3.705 186.295 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 190.285 3.705 190.855 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 202.065 3.705 202.635 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 197.695 3.705 198.265 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 194.845 3.705 195.415 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 207.005 4.465 207.575 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 207.765 4.465 208.335 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 208.145 3.705 208.715 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 198.455 3.705 199.025 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 185.345 4.465 185.915 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 190.665 4.465 191.235 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 193.895 3.705 194.465 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 191.045 3.705 191.615 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 188.955 3.705 189.525 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 186.485 3.705 187.055 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 184.965 3.705 185.535 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 13.015 208.525 13.585 209.095 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 14.155 208.525 14.725 209.095 ;
  END
 END i18
 PIN i19
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 13.015 195.225 13.585 195.795 ;
  END
 END i19
 PIN i20
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 14.155 195.225 14.725 195.795 ;
  END
 END i20
 PIN i21
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 401.755 26.885 402.325 ;
  END
 END i21
 PIN i22
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 385.415 26.885 385.985 ;
  END
 END i22
 PIN i23
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 220.115 26.885 220.685 ;
  END
 END i23
 PIN i24
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 172.235 26.885 172.805 ;
  END
 END i24
 PIN i25
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 155.895 26.885 156.465 ;
  END
 END i25
 PIN i26
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 139.555 26.885 140.125 ;
  END
 END i26
 PIN i27
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 123.215 26.885 123.785 ;
  END
 END i27
 PIN i28
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 106.875 26.885 107.445 ;
  END
 END i28
 PIN i29
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 72.295 26.885 72.865 ;
  END
 END i29
 PIN i30
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 55.955 26.885 56.525 ;
  END
 END i30
 PIN i31
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 39.615 26.885 40.185 ;
  END
 END i31
 PIN i32
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 23.275 26.885 23.845 ;
  END
 END i32
 PIN i33
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 369.075 26.885 369.645 ;
  END
 END i33
 PIN i34
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 6.935 26.885 7.505 ;
  END
 END i34
 PIN i35
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 352.735 26.885 353.305 ;
  END
 END i35
 PIN i36
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 336.395 26.885 336.965 ;
  END
 END i36
 PIN i37
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 320.055 26.885 320.625 ;
  END
 END i37
 PIN i38
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 285.475 26.885 286.045 ;
  END
 END i38
 PIN i39
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 269.135 26.885 269.705 ;
  END
 END i39
 PIN i40
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 252.795 26.885 253.365 ;
  END
 END i40
 PIN i41
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 236.455 26.885 237.025 ;
  END
 END i41
 PIN i42
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 334.115 27.645 334.685 ;
  END
 END i42
 PIN i43
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 330.125 26.885 330.695 ;
  END
 END i43
 PIN i44
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 325.945 26.885 326.515 ;
  END
 END i44
 PIN i45
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 346.465 26.885 347.035 ;
  END
 END i45
 PIN i46
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 342.285 26.885 342.855 ;
  END
 END i46
 PIN i47
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 266.855 27.645 267.425 ;
  END
 END i47
 PIN i48
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 262.865 26.885 263.435 ;
  END
 END i48
 PIN i49
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 258.685 26.885 259.255 ;
  END
 END i49
 PIN i50
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 254.695 26.885 255.265 ;
  END
 END i50
 PIN i51
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 250.515 27.645 251.085 ;
  END
 END i51
 PIN i52
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 125.495 27.645 126.065 ;
  END
 END i52
 PIN i53
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 129.485 26.885 130.055 ;
  END
 END i53
 PIN i54
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 133.665 26.885 134.235 ;
  END
 END i54
 PIN i55
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 137.655 26.885 138.225 ;
  END
 END i55
 PIN i56
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 141.835 27.645 142.405 ;
  END
 END i56
 PIN i57
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 58.235 27.645 58.805 ;
  END
 END i57
 PIN i58
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 62.225 26.885 62.795 ;
  END
 END i58
 PIN i59
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 66.405 26.885 66.975 ;
  END
 END i59
 PIN i60
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 45.885 26.885 46.455 ;
  END
 END i60
 PIN i61
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 50.065 26.885 50.635 ;
  END
 END i61
 PIN i62
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 338.295 26.885 338.865 ;
  END
 END i62
 PIN i63
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 271.035 26.885 271.605 ;
  END
 END i63
 PIN i64
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 121.315 26.885 121.885 ;
  END
 END i64
 PIN i65
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 54.055 26.885 54.625 ;
  END
 END i65
 PIN i66
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 18.335 208.525 18.905 209.095 ;
  END
 END i66
 PIN i67
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 18.335 195.225 18.905 195.795 ;
  END
 END i67
 PIN i68
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 401.185 27.645 401.755 ;
  END
 END i68
 PIN i69
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 384.845 27.645 385.415 ;
  END
 END i69
 PIN i70
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 219.545 27.645 220.115 ;
  END
 END i70
 PIN i71
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 172.805 27.645 173.375 ;
  END
 END i71
 PIN i72
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 156.465 27.645 157.035 ;
  END
 END i72
 PIN i73
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 140.125 27.645 140.695 ;
  END
 END i73
 PIN i74
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 123.785 27.645 124.355 ;
  END
 END i74
 PIN i75
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 107.445 27.645 108.015 ;
  END
 END i75
 PIN i76
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 72.865 27.645 73.435 ;
  END
 END i76
 PIN i77
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 56.525 27.645 57.095 ;
  END
 END i77
 PIN i78
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 40.185 27.645 40.755 ;
  END
 END i78
 PIN i79
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 23.845 27.645 24.415 ;
  END
 END i79
 PIN i80
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 368.505 27.645 369.075 ;
  END
 END i80
 PIN i81
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 7.505 27.645 8.075 ;
  END
 END i81
 PIN i82
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 352.165 27.645 352.735 ;
  END
 END i82
 PIN i83
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 335.825 27.645 336.395 ;
  END
 END i83
 PIN i84
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 319.485 27.645 320.055 ;
  END
 END i84
 PIN i85
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 284.905 27.645 285.475 ;
  END
 END i85
 PIN i86
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 268.565 27.645 269.135 ;
  END
 END i86
 PIN i87
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 252.225 27.645 252.795 ;
  END
 END i87
 PIN i88
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 235.885 27.645 236.455 ;
  END
 END i88
 PIN i89
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 200.925 3.705 201.495 ;
  END
 END i89
 PIN i90
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 200.545 4.465 201.115 ;
  END
 END i90
 PIN i91
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 400.615 28.405 401.185 ;
  END
 END i91
 PIN i92
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 384.275 28.405 384.845 ;
  END
 END i92
 PIN i93
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 218.975 28.405 219.545 ;
  END
 END i93
 PIN i94
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 173.375 28.405 173.945 ;
  END
 END i94
 PIN i95
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 157.035 28.405 157.605 ;
  END
 END i95
 PIN i96
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 140.695 28.405 141.265 ;
  END
 END i96
 PIN i97
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 124.355 28.405 124.925 ;
  END
 END i97
 PIN i98
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 108.015 28.405 108.585 ;
  END
 END i98
 PIN i99
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 73.435 28.405 74.005 ;
  END
 END i99
 PIN i100
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 57.095 28.405 57.665 ;
  END
 END i100
 PIN i101
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 40.755 28.405 41.325 ;
  END
 END i101
 PIN i102
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 24.415 28.405 24.985 ;
  END
 END i102
 PIN i103
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 367.935 28.405 368.505 ;
  END
 END i103
 PIN i104
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 8.075 28.405 8.645 ;
  END
 END i104
 PIN i105
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 351.595 28.405 352.165 ;
  END
 END i105
 PIN i106
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 335.255 28.405 335.825 ;
  END
 END i106
 PIN i107
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 318.915 28.405 319.485 ;
  END
 END i107
 PIN i108
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 284.335 28.405 284.905 ;
  END
 END i108
 PIN i109
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 267.995 28.405 268.565 ;
  END
 END i109
 PIN i110
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 251.655 28.405 252.225 ;
  END
 END i110
 PIN i111
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 235.315 28.405 235.885 ;
  END
 END i111
 PIN i112
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 4.275 208.525 4.845 209.095 ;
  END
 END i112
 PIN i113
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 5.415 208.525 5.985 209.095 ;
  END
 END i113
 PIN i114
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 7.315 208.525 7.885 209.095 ;
  END
 END i114
 PIN i115
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 8.835 208.525 9.405 209.095 ;
  END
 END i115
 PIN i116
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 208.525 10.925 209.095 ;
  END
 END i116
 PIN i117
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 11.875 208.525 12.445 209.095 ;
  END
 END i117
 PIN i118
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 4.275 195.225 4.845 195.795 ;
  END
 END i118
 PIN i119
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 5.415 195.225 5.985 195.795 ;
  END
 END i119
 PIN i120
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 7.315 195.225 7.885 195.795 ;
  END
 END i120
 PIN i121
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 8.835 195.225 9.405 195.795 ;
  END
 END i121
 PIN i122
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 195.225 10.925 195.795 ;
  END
 END i122
 PIN i123
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 11.875 195.225 12.445 195.795 ;
  END
 END i123
 OBS
  LAYER metal1 ;
   RECT 23.18 0.0 508.44 1.71 ;
   RECT 23.18 1.71 508.44 3.42 ;
   RECT 23.18 3.42 508.44 5.13 ;
   RECT 23.18 5.13 508.44 6.84 ;
   RECT 23.18 6.84 508.44 8.55 ;
   RECT 23.18 8.55 508.44 10.26 ;
   RECT 23.18 10.26 508.44 11.97 ;
   RECT 23.18 11.97 508.44 13.68 ;
   RECT 23.18 13.68 508.44 15.39 ;
   RECT 23.18 15.39 508.44 17.1 ;
   RECT 23.18 17.1 508.44 18.81 ;
   RECT 23.18 18.81 508.44 20.52 ;
   RECT 23.18 20.52 508.44 22.23 ;
   RECT 23.18 22.23 508.44 23.94 ;
   RECT 23.18 23.94 508.44 25.65 ;
   RECT 23.18 25.65 508.44 27.36 ;
   RECT 23.18 27.36 508.44 29.07 ;
   RECT 23.18 29.07 508.44 30.78 ;
   RECT 23.18 30.78 508.44 32.49 ;
   RECT 23.18 32.49 508.44 34.2 ;
   RECT 23.18 34.2 508.44 35.91 ;
   RECT 23.18 35.91 508.44 37.62 ;
   RECT 23.18 37.62 508.44 39.33 ;
   RECT 23.18 39.33 508.44 41.04 ;
   RECT 23.18 41.04 508.44 42.75 ;
   RECT 23.18 42.75 508.44 44.46 ;
   RECT 23.18 44.46 508.44 46.17 ;
   RECT 23.18 46.17 508.44 47.88 ;
   RECT 23.18 47.88 508.44 49.59 ;
   RECT 23.18 49.59 508.44 51.3 ;
   RECT 23.18 51.3 508.44 53.01 ;
   RECT 23.18 53.01 508.44 54.72 ;
   RECT 23.18 54.72 508.44 56.43 ;
   RECT 23.18 56.43 508.44 58.14 ;
   RECT 23.18 58.14 508.44 59.85 ;
   RECT 23.18 59.85 508.44 61.56 ;
   RECT 23.18 61.56 508.44 63.27 ;
   RECT 23.18 63.27 508.44 64.98 ;
   RECT 23.18 64.98 508.44 66.69 ;
   RECT 23.18 66.69 508.44 68.4 ;
   RECT 23.18 68.4 508.44 70.11 ;
   RECT 23.18 70.11 508.44 71.82 ;
   RECT 23.18 71.82 508.44 73.53 ;
   RECT 23.18 73.53 508.44 75.24 ;
   RECT 23.18 75.24 508.44 76.95 ;
   RECT 23.18 76.95 508.44 78.66 ;
   RECT 23.18 78.66 508.44 80.37 ;
   RECT 23.18 80.37 508.44 82.08 ;
   RECT 23.18 82.08 508.44 83.79 ;
   RECT 23.18 83.79 508.44 85.5 ;
   RECT 23.18 85.5 508.44 87.21 ;
   RECT 23.18 87.21 508.44 88.92 ;
   RECT 23.18 88.92 508.44 90.63 ;
   RECT 23.18 90.63 508.44 92.34 ;
   RECT 23.18 92.34 508.44 94.05 ;
   RECT 23.18 94.05 508.44 95.76 ;
   RECT 23.18 95.76 508.44 97.47 ;
   RECT 23.18 97.47 508.44 99.18 ;
   RECT 23.18 99.18 508.44 100.89 ;
   RECT 23.18 100.89 508.44 102.6 ;
   RECT 23.18 102.6 508.44 104.31 ;
   RECT 23.18 104.31 508.44 106.02 ;
   RECT 23.18 106.02 508.44 107.73 ;
   RECT 23.18 107.73 508.44 109.44 ;
   RECT 23.18 109.44 508.44 111.15 ;
   RECT 23.18 111.15 508.44 112.86 ;
   RECT 23.18 112.86 508.44 114.57 ;
   RECT 23.18 114.57 508.44 116.28 ;
   RECT 23.18 116.28 508.44 117.99 ;
   RECT 23.18 117.99 508.44 119.7 ;
   RECT 23.18 119.7 508.44 121.41 ;
   RECT 23.18 121.41 508.44 123.12 ;
   RECT 23.18 123.12 508.44 124.83 ;
   RECT 23.18 124.83 508.44 126.54 ;
   RECT 23.18 126.54 508.44 128.25 ;
   RECT 23.18 128.25 508.44 129.96 ;
   RECT 23.18 129.96 508.44 131.67 ;
   RECT 23.18 131.67 508.44 133.38 ;
   RECT 23.18 133.38 508.44 135.09 ;
   RECT 23.18 135.09 508.44 136.8 ;
   RECT 23.18 136.8 508.44 138.51 ;
   RECT 23.18 138.51 508.44 140.22 ;
   RECT 23.18 140.22 508.44 141.93 ;
   RECT 23.18 141.93 508.44 143.64 ;
   RECT 23.18 143.64 508.44 145.35 ;
   RECT 23.18 145.35 508.44 147.06 ;
   RECT 23.18 147.06 508.44 148.77 ;
   RECT 23.18 148.77 508.44 150.48 ;
   RECT 23.18 150.48 508.44 152.19 ;
   RECT 23.18 152.19 508.44 153.9 ;
   RECT 23.18 153.9 508.44 155.61 ;
   RECT 23.18 155.61 508.44 157.32 ;
   RECT 23.18 157.32 508.44 159.03 ;
   RECT 23.18 159.03 508.44 160.74 ;
   RECT 23.18 160.74 508.44 162.45 ;
   RECT 23.18 162.45 508.44 164.16 ;
   RECT 23.18 164.16 508.44 165.87 ;
   RECT 23.18 165.87 508.44 167.58 ;
   RECT 23.18 167.58 508.44 169.29 ;
   RECT 23.18 169.29 508.44 171.0 ;
   RECT 23.18 171.0 508.44 172.71 ;
   RECT 23.18 172.71 508.44 174.42 ;
   RECT 23.18 174.42 508.44 176.13 ;
   RECT 23.18 176.13 508.44 177.84 ;
   RECT 23.18 177.84 508.44 179.55 ;
   RECT 23.18 179.55 508.44 181.26 ;
   RECT 23.18 181.26 508.44 182.97 ;
   RECT 0.0 182.97 508.44 184.68 ;
   RECT 0.0 184.68 508.44 186.39 ;
   RECT 0.0 186.39 508.44 188.1 ;
   RECT 0.0 188.1 508.44 189.81 ;
   RECT 0.0 189.81 508.44 191.52 ;
   RECT 0.0 191.52 508.44 193.23 ;
   RECT 0.0 193.23 508.44 194.94 ;
   RECT 0.0 194.94 508.44 196.65 ;
   RECT 0.0 196.65 508.44 198.36 ;
   RECT 0.0 198.36 508.44 200.07 ;
   RECT 0.0 200.07 508.44 201.78 ;
   RECT 0.0 201.78 508.44 203.49 ;
   RECT 0.0 203.49 508.44 205.2 ;
   RECT 0.0 205.2 508.44 206.91 ;
   RECT 0.0 206.91 508.44 208.62 ;
   RECT 0.0 208.62 508.44 210.33 ;
   RECT 0.0 210.33 508.44 212.04 ;
   RECT 23.18 212.04 508.44 213.75 ;
   RECT 23.18 213.75 508.44 215.46 ;
   RECT 23.18 215.46 508.44 217.17 ;
   RECT 23.18 217.17 508.44 218.88 ;
   RECT 23.18 218.88 508.44 220.59 ;
   RECT 23.18 220.59 508.44 222.3 ;
   RECT 23.18 222.3 508.44 224.01 ;
   RECT 23.18 224.01 508.44 225.72 ;
   RECT 23.18 225.72 508.44 227.43 ;
   RECT 23.18 227.43 508.44 229.14 ;
   RECT 23.18 229.14 508.44 230.85 ;
   RECT 23.18 230.85 508.44 232.56 ;
   RECT 23.18 232.56 508.44 234.27 ;
   RECT 23.18 234.27 508.44 235.98 ;
   RECT 23.18 235.98 508.44 237.69 ;
   RECT 23.18 237.69 508.44 239.4 ;
   RECT 23.18 239.4 508.44 241.11 ;
   RECT 23.18 241.11 508.44 242.82 ;
   RECT 23.18 242.82 508.44 244.53 ;
   RECT 23.18 244.53 508.44 246.24 ;
   RECT 23.18 246.24 508.44 247.95 ;
   RECT 23.18 247.95 508.44 249.66 ;
   RECT 23.18 249.66 508.44 251.37 ;
   RECT 23.18 251.37 508.44 253.08 ;
   RECT 23.18 253.08 508.44 254.79 ;
   RECT 23.18 254.79 508.44 256.5 ;
   RECT 23.18 256.5 508.44 258.21 ;
   RECT 23.18 258.21 508.44 259.92 ;
   RECT 23.18 259.92 508.44 261.63 ;
   RECT 23.18 261.63 508.44 263.34 ;
   RECT 23.18 263.34 508.44 265.05 ;
   RECT 23.18 265.05 508.44 266.76 ;
   RECT 23.18 266.76 508.44 268.47 ;
   RECT 23.18 268.47 508.44 270.18 ;
   RECT 23.18 270.18 508.44 271.89 ;
   RECT 23.18 271.89 508.44 273.6 ;
   RECT 23.18 273.6 508.44 275.31 ;
   RECT 23.18 275.31 508.44 277.02 ;
   RECT 23.18 277.02 508.44 278.73 ;
   RECT 23.18 278.73 508.44 280.44 ;
   RECT 23.18 280.44 508.44 282.15 ;
   RECT 23.18 282.15 508.44 283.86 ;
   RECT 23.18 283.86 508.44 285.57 ;
   RECT 23.18 285.57 508.44 287.28 ;
   RECT 23.18 287.28 508.44 288.99 ;
   RECT 23.18 288.99 508.44 290.7 ;
   RECT 23.18 290.7 508.44 292.41 ;
   RECT 23.18 292.41 508.44 294.12 ;
   RECT 23.18 294.12 508.44 295.83 ;
   RECT 23.18 295.83 508.44 297.54 ;
   RECT 23.18 297.54 508.44 299.25 ;
   RECT 23.18 299.25 508.44 300.96 ;
   RECT 23.18 300.96 508.44 302.67 ;
   RECT 23.18 302.67 508.44 304.38 ;
   RECT 23.18 304.38 508.44 306.09 ;
   RECT 23.18 306.09 508.44 307.8 ;
   RECT 23.18 307.8 508.44 309.51 ;
   RECT 23.18 309.51 508.44 311.22 ;
   RECT 23.18 311.22 508.44 312.93 ;
   RECT 23.18 312.93 508.44 314.64 ;
   RECT 23.18 314.64 508.44 316.35 ;
   RECT 23.18 316.35 508.44 318.06 ;
   RECT 23.18 318.06 508.44 319.77 ;
   RECT 23.18 319.77 508.44 321.48 ;
   RECT 23.18 321.48 508.44 323.19 ;
   RECT 23.18 323.19 508.44 324.9 ;
   RECT 23.18 324.9 508.44 326.61 ;
   RECT 23.18 326.61 508.44 328.32 ;
   RECT 23.18 328.32 508.44 330.03 ;
   RECT 23.18 330.03 508.44 331.74 ;
   RECT 23.18 331.74 508.44 333.45 ;
   RECT 23.18 333.45 508.44 335.16 ;
   RECT 23.18 335.16 508.44 336.87 ;
   RECT 23.18 336.87 508.44 338.58 ;
   RECT 23.18 338.58 508.44 340.29 ;
   RECT 23.18 340.29 508.44 342.0 ;
   RECT 23.18 342.0 508.44 343.71 ;
   RECT 23.18 343.71 508.44 345.42 ;
   RECT 23.18 345.42 508.44 347.13 ;
   RECT 23.18 347.13 508.44 348.84 ;
   RECT 23.18 348.84 508.44 350.55 ;
   RECT 23.18 350.55 508.44 352.26 ;
   RECT 23.18 352.26 508.44 353.97 ;
   RECT 23.18 353.97 508.44 355.68 ;
   RECT 23.18 355.68 508.44 357.39 ;
   RECT 23.18 357.39 508.44 359.1 ;
   RECT 23.18 359.1 508.44 360.81 ;
   RECT 23.18 360.81 508.44 362.52 ;
   RECT 23.18 362.52 508.44 364.23 ;
   RECT 23.18 364.23 508.44 365.94 ;
   RECT 23.18 365.94 508.44 367.65 ;
   RECT 23.18 367.65 508.44 369.36 ;
   RECT 23.18 369.36 508.44 371.07 ;
   RECT 23.18 371.07 508.44 372.78 ;
   RECT 23.18 372.78 508.44 374.49 ;
   RECT 23.18 374.49 508.44 376.2 ;
   RECT 23.18 376.2 508.44 377.91 ;
   RECT 23.18 377.91 508.44 379.62 ;
   RECT 23.18 379.62 508.44 381.33 ;
   RECT 23.18 381.33 508.44 383.04 ;
   RECT 23.18 383.04 508.44 384.75 ;
   RECT 23.18 384.75 508.44 386.46 ;
   RECT 23.18 386.46 508.44 388.17 ;
   RECT 23.18 388.17 508.44 389.88 ;
   RECT 23.18 389.88 508.44 391.59 ;
   RECT 23.18 391.59 508.44 393.3 ;
   RECT 23.18 393.3 508.44 395.01 ;
   RECT 23.18 395.01 508.44 396.72 ;
   RECT 23.18 396.72 508.44 398.43 ;
   RECT 23.18 398.43 508.44 400.14 ;
   RECT 23.18 400.14 508.44 401.85 ;
   RECT 23.18 401.85 508.44 403.56 ;
   RECT 23.18 403.56 508.44 405.27 ;
   RECT 23.18 405.27 508.44 406.98 ;
   RECT 23.18 406.98 508.44 408.69 ;
   RECT 23.18 408.69 508.44 410.4 ;
  LAYER via1 ;
   RECT 23.18 0.0 508.44 1.71 ;
   RECT 23.18 1.71 508.44 3.42 ;
   RECT 23.18 3.42 508.44 5.13 ;
   RECT 23.18 5.13 508.44 6.84 ;
   RECT 23.18 6.84 508.44 8.55 ;
   RECT 23.18 8.55 508.44 10.26 ;
   RECT 23.18 10.26 508.44 11.97 ;
   RECT 23.18 11.97 508.44 13.68 ;
   RECT 23.18 13.68 508.44 15.39 ;
   RECT 23.18 15.39 508.44 17.1 ;
   RECT 23.18 17.1 508.44 18.81 ;
   RECT 23.18 18.81 508.44 20.52 ;
   RECT 23.18 20.52 508.44 22.23 ;
   RECT 23.18 22.23 508.44 23.94 ;
   RECT 23.18 23.94 508.44 25.65 ;
   RECT 23.18 25.65 508.44 27.36 ;
   RECT 23.18 27.36 508.44 29.07 ;
   RECT 23.18 29.07 508.44 30.78 ;
   RECT 23.18 30.78 508.44 32.49 ;
   RECT 23.18 32.49 508.44 34.2 ;
   RECT 23.18 34.2 508.44 35.91 ;
   RECT 23.18 35.91 508.44 37.62 ;
   RECT 23.18 37.62 508.44 39.33 ;
   RECT 23.18 39.33 508.44 41.04 ;
   RECT 23.18 41.04 508.44 42.75 ;
   RECT 23.18 42.75 508.44 44.46 ;
   RECT 23.18 44.46 508.44 46.17 ;
   RECT 23.18 46.17 508.44 47.88 ;
   RECT 23.18 47.88 508.44 49.59 ;
   RECT 23.18 49.59 508.44 51.3 ;
   RECT 23.18 51.3 508.44 53.01 ;
   RECT 23.18 53.01 508.44 54.72 ;
   RECT 23.18 54.72 508.44 56.43 ;
   RECT 23.18 56.43 508.44 58.14 ;
   RECT 23.18 58.14 508.44 59.85 ;
   RECT 23.18 59.85 508.44 61.56 ;
   RECT 23.18 61.56 508.44 63.27 ;
   RECT 23.18 63.27 508.44 64.98 ;
   RECT 23.18 64.98 508.44 66.69 ;
   RECT 23.18 66.69 508.44 68.4 ;
   RECT 23.18 68.4 508.44 70.11 ;
   RECT 23.18 70.11 508.44 71.82 ;
   RECT 23.18 71.82 508.44 73.53 ;
   RECT 23.18 73.53 508.44 75.24 ;
   RECT 23.18 75.24 508.44 76.95 ;
   RECT 23.18 76.95 508.44 78.66 ;
   RECT 23.18 78.66 508.44 80.37 ;
   RECT 23.18 80.37 508.44 82.08 ;
   RECT 23.18 82.08 508.44 83.79 ;
   RECT 23.18 83.79 508.44 85.5 ;
   RECT 23.18 85.5 508.44 87.21 ;
   RECT 23.18 87.21 508.44 88.92 ;
   RECT 23.18 88.92 508.44 90.63 ;
   RECT 23.18 90.63 508.44 92.34 ;
   RECT 23.18 92.34 508.44 94.05 ;
   RECT 23.18 94.05 508.44 95.76 ;
   RECT 23.18 95.76 508.44 97.47 ;
   RECT 23.18 97.47 508.44 99.18 ;
   RECT 23.18 99.18 508.44 100.89 ;
   RECT 23.18 100.89 508.44 102.6 ;
   RECT 23.18 102.6 508.44 104.31 ;
   RECT 23.18 104.31 508.44 106.02 ;
   RECT 23.18 106.02 508.44 107.73 ;
   RECT 23.18 107.73 508.44 109.44 ;
   RECT 23.18 109.44 508.44 111.15 ;
   RECT 23.18 111.15 508.44 112.86 ;
   RECT 23.18 112.86 508.44 114.57 ;
   RECT 23.18 114.57 508.44 116.28 ;
   RECT 23.18 116.28 508.44 117.99 ;
   RECT 23.18 117.99 508.44 119.7 ;
   RECT 23.18 119.7 508.44 121.41 ;
   RECT 23.18 121.41 508.44 123.12 ;
   RECT 23.18 123.12 508.44 124.83 ;
   RECT 23.18 124.83 508.44 126.54 ;
   RECT 23.18 126.54 508.44 128.25 ;
   RECT 23.18 128.25 508.44 129.96 ;
   RECT 23.18 129.96 508.44 131.67 ;
   RECT 23.18 131.67 508.44 133.38 ;
   RECT 23.18 133.38 508.44 135.09 ;
   RECT 23.18 135.09 508.44 136.8 ;
   RECT 23.18 136.8 508.44 138.51 ;
   RECT 23.18 138.51 508.44 140.22 ;
   RECT 23.18 140.22 508.44 141.93 ;
   RECT 23.18 141.93 508.44 143.64 ;
   RECT 23.18 143.64 508.44 145.35 ;
   RECT 23.18 145.35 508.44 147.06 ;
   RECT 23.18 147.06 508.44 148.77 ;
   RECT 23.18 148.77 508.44 150.48 ;
   RECT 23.18 150.48 508.44 152.19 ;
   RECT 23.18 152.19 508.44 153.9 ;
   RECT 23.18 153.9 508.44 155.61 ;
   RECT 23.18 155.61 508.44 157.32 ;
   RECT 23.18 157.32 508.44 159.03 ;
   RECT 23.18 159.03 508.44 160.74 ;
   RECT 23.18 160.74 508.44 162.45 ;
   RECT 23.18 162.45 508.44 164.16 ;
   RECT 23.18 164.16 508.44 165.87 ;
   RECT 23.18 165.87 508.44 167.58 ;
   RECT 23.18 167.58 508.44 169.29 ;
   RECT 23.18 169.29 508.44 171.0 ;
   RECT 23.18 171.0 508.44 172.71 ;
   RECT 23.18 172.71 508.44 174.42 ;
   RECT 23.18 174.42 508.44 176.13 ;
   RECT 23.18 176.13 508.44 177.84 ;
   RECT 23.18 177.84 508.44 179.55 ;
   RECT 23.18 179.55 508.44 181.26 ;
   RECT 23.18 181.26 508.44 182.97 ;
   RECT 0.0 182.97 508.44 184.68 ;
   RECT 0.0 184.68 508.44 186.39 ;
   RECT 0.0 186.39 508.44 188.1 ;
   RECT 0.0 188.1 508.44 189.81 ;
   RECT 0.0 189.81 508.44 191.52 ;
   RECT 0.0 191.52 508.44 193.23 ;
   RECT 0.0 193.23 508.44 194.94 ;
   RECT 0.0 194.94 508.44 196.65 ;
   RECT 0.0 196.65 508.44 198.36 ;
   RECT 0.0 198.36 508.44 200.07 ;
   RECT 0.0 200.07 508.44 201.78 ;
   RECT 0.0 201.78 508.44 203.49 ;
   RECT 0.0 203.49 508.44 205.2 ;
   RECT 0.0 205.2 508.44 206.91 ;
   RECT 0.0 206.91 508.44 208.62 ;
   RECT 0.0 208.62 508.44 210.33 ;
   RECT 0.0 210.33 508.44 212.04 ;
   RECT 23.18 212.04 508.44 213.75 ;
   RECT 23.18 213.75 508.44 215.46 ;
   RECT 23.18 215.46 508.44 217.17 ;
   RECT 23.18 217.17 508.44 218.88 ;
   RECT 23.18 218.88 508.44 220.59 ;
   RECT 23.18 220.59 508.44 222.3 ;
   RECT 23.18 222.3 508.44 224.01 ;
   RECT 23.18 224.01 508.44 225.72 ;
   RECT 23.18 225.72 508.44 227.43 ;
   RECT 23.18 227.43 508.44 229.14 ;
   RECT 23.18 229.14 508.44 230.85 ;
   RECT 23.18 230.85 508.44 232.56 ;
   RECT 23.18 232.56 508.44 234.27 ;
   RECT 23.18 234.27 508.44 235.98 ;
   RECT 23.18 235.98 508.44 237.69 ;
   RECT 23.18 237.69 508.44 239.4 ;
   RECT 23.18 239.4 508.44 241.11 ;
   RECT 23.18 241.11 508.44 242.82 ;
   RECT 23.18 242.82 508.44 244.53 ;
   RECT 23.18 244.53 508.44 246.24 ;
   RECT 23.18 246.24 508.44 247.95 ;
   RECT 23.18 247.95 508.44 249.66 ;
   RECT 23.18 249.66 508.44 251.37 ;
   RECT 23.18 251.37 508.44 253.08 ;
   RECT 23.18 253.08 508.44 254.79 ;
   RECT 23.18 254.79 508.44 256.5 ;
   RECT 23.18 256.5 508.44 258.21 ;
   RECT 23.18 258.21 508.44 259.92 ;
   RECT 23.18 259.92 508.44 261.63 ;
   RECT 23.18 261.63 508.44 263.34 ;
   RECT 23.18 263.34 508.44 265.05 ;
   RECT 23.18 265.05 508.44 266.76 ;
   RECT 23.18 266.76 508.44 268.47 ;
   RECT 23.18 268.47 508.44 270.18 ;
   RECT 23.18 270.18 508.44 271.89 ;
   RECT 23.18 271.89 508.44 273.6 ;
   RECT 23.18 273.6 508.44 275.31 ;
   RECT 23.18 275.31 508.44 277.02 ;
   RECT 23.18 277.02 508.44 278.73 ;
   RECT 23.18 278.73 508.44 280.44 ;
   RECT 23.18 280.44 508.44 282.15 ;
   RECT 23.18 282.15 508.44 283.86 ;
   RECT 23.18 283.86 508.44 285.57 ;
   RECT 23.18 285.57 508.44 287.28 ;
   RECT 23.18 287.28 508.44 288.99 ;
   RECT 23.18 288.99 508.44 290.7 ;
   RECT 23.18 290.7 508.44 292.41 ;
   RECT 23.18 292.41 508.44 294.12 ;
   RECT 23.18 294.12 508.44 295.83 ;
   RECT 23.18 295.83 508.44 297.54 ;
   RECT 23.18 297.54 508.44 299.25 ;
   RECT 23.18 299.25 508.44 300.96 ;
   RECT 23.18 300.96 508.44 302.67 ;
   RECT 23.18 302.67 508.44 304.38 ;
   RECT 23.18 304.38 508.44 306.09 ;
   RECT 23.18 306.09 508.44 307.8 ;
   RECT 23.18 307.8 508.44 309.51 ;
   RECT 23.18 309.51 508.44 311.22 ;
   RECT 23.18 311.22 508.44 312.93 ;
   RECT 23.18 312.93 508.44 314.64 ;
   RECT 23.18 314.64 508.44 316.35 ;
   RECT 23.18 316.35 508.44 318.06 ;
   RECT 23.18 318.06 508.44 319.77 ;
   RECT 23.18 319.77 508.44 321.48 ;
   RECT 23.18 321.48 508.44 323.19 ;
   RECT 23.18 323.19 508.44 324.9 ;
   RECT 23.18 324.9 508.44 326.61 ;
   RECT 23.18 326.61 508.44 328.32 ;
   RECT 23.18 328.32 508.44 330.03 ;
   RECT 23.18 330.03 508.44 331.74 ;
   RECT 23.18 331.74 508.44 333.45 ;
   RECT 23.18 333.45 508.44 335.16 ;
   RECT 23.18 335.16 508.44 336.87 ;
   RECT 23.18 336.87 508.44 338.58 ;
   RECT 23.18 338.58 508.44 340.29 ;
   RECT 23.18 340.29 508.44 342.0 ;
   RECT 23.18 342.0 508.44 343.71 ;
   RECT 23.18 343.71 508.44 345.42 ;
   RECT 23.18 345.42 508.44 347.13 ;
   RECT 23.18 347.13 508.44 348.84 ;
   RECT 23.18 348.84 508.44 350.55 ;
   RECT 23.18 350.55 508.44 352.26 ;
   RECT 23.18 352.26 508.44 353.97 ;
   RECT 23.18 353.97 508.44 355.68 ;
   RECT 23.18 355.68 508.44 357.39 ;
   RECT 23.18 357.39 508.44 359.1 ;
   RECT 23.18 359.1 508.44 360.81 ;
   RECT 23.18 360.81 508.44 362.52 ;
   RECT 23.18 362.52 508.44 364.23 ;
   RECT 23.18 364.23 508.44 365.94 ;
   RECT 23.18 365.94 508.44 367.65 ;
   RECT 23.18 367.65 508.44 369.36 ;
   RECT 23.18 369.36 508.44 371.07 ;
   RECT 23.18 371.07 508.44 372.78 ;
   RECT 23.18 372.78 508.44 374.49 ;
   RECT 23.18 374.49 508.44 376.2 ;
   RECT 23.18 376.2 508.44 377.91 ;
   RECT 23.18 377.91 508.44 379.62 ;
   RECT 23.18 379.62 508.44 381.33 ;
   RECT 23.18 381.33 508.44 383.04 ;
   RECT 23.18 383.04 508.44 384.75 ;
   RECT 23.18 384.75 508.44 386.46 ;
   RECT 23.18 386.46 508.44 388.17 ;
   RECT 23.18 388.17 508.44 389.88 ;
   RECT 23.18 389.88 508.44 391.59 ;
   RECT 23.18 391.59 508.44 393.3 ;
   RECT 23.18 393.3 508.44 395.01 ;
   RECT 23.18 395.01 508.44 396.72 ;
   RECT 23.18 396.72 508.44 398.43 ;
   RECT 23.18 398.43 508.44 400.14 ;
   RECT 23.18 400.14 508.44 401.85 ;
   RECT 23.18 401.85 508.44 403.56 ;
   RECT 23.18 403.56 508.44 405.27 ;
   RECT 23.18 405.27 508.44 406.98 ;
   RECT 23.18 406.98 508.44 408.69 ;
   RECT 23.18 408.69 508.44 410.4 ;
  LAYER metal2 ;
   RECT 23.18 0.0 508.44 1.71 ;
   RECT 23.18 1.71 508.44 3.42 ;
   RECT 23.18 3.42 508.44 5.13 ;
   RECT 23.18 5.13 508.44 6.84 ;
   RECT 23.18 6.84 508.44 8.55 ;
   RECT 23.18 8.55 508.44 10.26 ;
   RECT 23.18 10.26 508.44 11.97 ;
   RECT 23.18 11.97 508.44 13.68 ;
   RECT 23.18 13.68 508.44 15.39 ;
   RECT 23.18 15.39 508.44 17.1 ;
   RECT 23.18 17.1 508.44 18.81 ;
   RECT 23.18 18.81 508.44 20.52 ;
   RECT 23.18 20.52 508.44 22.23 ;
   RECT 23.18 22.23 508.44 23.94 ;
   RECT 23.18 23.94 508.44 25.65 ;
   RECT 23.18 25.65 508.44 27.36 ;
   RECT 23.18 27.36 508.44 29.07 ;
   RECT 23.18 29.07 508.44 30.78 ;
   RECT 23.18 30.78 508.44 32.49 ;
   RECT 23.18 32.49 508.44 34.2 ;
   RECT 23.18 34.2 508.44 35.91 ;
   RECT 23.18 35.91 508.44 37.62 ;
   RECT 23.18 37.62 508.44 39.33 ;
   RECT 23.18 39.33 508.44 41.04 ;
   RECT 23.18 41.04 508.44 42.75 ;
   RECT 23.18 42.75 508.44 44.46 ;
   RECT 23.18 44.46 508.44 46.17 ;
   RECT 23.18 46.17 508.44 47.88 ;
   RECT 23.18 47.88 508.44 49.59 ;
   RECT 23.18 49.59 508.44 51.3 ;
   RECT 23.18 51.3 508.44 53.01 ;
   RECT 23.18 53.01 508.44 54.72 ;
   RECT 23.18 54.72 508.44 56.43 ;
   RECT 23.18 56.43 508.44 58.14 ;
   RECT 23.18 58.14 508.44 59.85 ;
   RECT 23.18 59.85 508.44 61.56 ;
   RECT 23.18 61.56 508.44 63.27 ;
   RECT 23.18 63.27 508.44 64.98 ;
   RECT 23.18 64.98 508.44 66.69 ;
   RECT 23.18 66.69 508.44 68.4 ;
   RECT 23.18 68.4 508.44 70.11 ;
   RECT 23.18 70.11 508.44 71.82 ;
   RECT 23.18 71.82 508.44 73.53 ;
   RECT 23.18 73.53 508.44 75.24 ;
   RECT 23.18 75.24 508.44 76.95 ;
   RECT 23.18 76.95 508.44 78.66 ;
   RECT 23.18 78.66 508.44 80.37 ;
   RECT 23.18 80.37 508.44 82.08 ;
   RECT 23.18 82.08 508.44 83.79 ;
   RECT 23.18 83.79 508.44 85.5 ;
   RECT 23.18 85.5 508.44 87.21 ;
   RECT 23.18 87.21 508.44 88.92 ;
   RECT 23.18 88.92 508.44 90.63 ;
   RECT 23.18 90.63 508.44 92.34 ;
   RECT 23.18 92.34 508.44 94.05 ;
   RECT 23.18 94.05 508.44 95.76 ;
   RECT 23.18 95.76 508.44 97.47 ;
   RECT 23.18 97.47 508.44 99.18 ;
   RECT 23.18 99.18 508.44 100.89 ;
   RECT 23.18 100.89 508.44 102.6 ;
   RECT 23.18 102.6 508.44 104.31 ;
   RECT 23.18 104.31 508.44 106.02 ;
   RECT 23.18 106.02 508.44 107.73 ;
   RECT 23.18 107.73 508.44 109.44 ;
   RECT 23.18 109.44 508.44 111.15 ;
   RECT 23.18 111.15 508.44 112.86 ;
   RECT 23.18 112.86 508.44 114.57 ;
   RECT 23.18 114.57 508.44 116.28 ;
   RECT 23.18 116.28 508.44 117.99 ;
   RECT 23.18 117.99 508.44 119.7 ;
   RECT 23.18 119.7 508.44 121.41 ;
   RECT 23.18 121.41 508.44 123.12 ;
   RECT 23.18 123.12 508.44 124.83 ;
   RECT 23.18 124.83 508.44 126.54 ;
   RECT 23.18 126.54 508.44 128.25 ;
   RECT 23.18 128.25 508.44 129.96 ;
   RECT 23.18 129.96 508.44 131.67 ;
   RECT 23.18 131.67 508.44 133.38 ;
   RECT 23.18 133.38 508.44 135.09 ;
   RECT 23.18 135.09 508.44 136.8 ;
   RECT 23.18 136.8 508.44 138.51 ;
   RECT 23.18 138.51 508.44 140.22 ;
   RECT 23.18 140.22 508.44 141.93 ;
   RECT 23.18 141.93 508.44 143.64 ;
   RECT 23.18 143.64 508.44 145.35 ;
   RECT 23.18 145.35 508.44 147.06 ;
   RECT 23.18 147.06 508.44 148.77 ;
   RECT 23.18 148.77 508.44 150.48 ;
   RECT 23.18 150.48 508.44 152.19 ;
   RECT 23.18 152.19 508.44 153.9 ;
   RECT 23.18 153.9 508.44 155.61 ;
   RECT 23.18 155.61 508.44 157.32 ;
   RECT 23.18 157.32 508.44 159.03 ;
   RECT 23.18 159.03 508.44 160.74 ;
   RECT 23.18 160.74 508.44 162.45 ;
   RECT 23.18 162.45 508.44 164.16 ;
   RECT 23.18 164.16 508.44 165.87 ;
   RECT 23.18 165.87 508.44 167.58 ;
   RECT 23.18 167.58 508.44 169.29 ;
   RECT 23.18 169.29 508.44 171.0 ;
   RECT 23.18 171.0 508.44 172.71 ;
   RECT 23.18 172.71 508.44 174.42 ;
   RECT 23.18 174.42 508.44 176.13 ;
   RECT 23.18 176.13 508.44 177.84 ;
   RECT 23.18 177.84 508.44 179.55 ;
   RECT 23.18 179.55 508.44 181.26 ;
   RECT 23.18 181.26 508.44 182.97 ;
   RECT 0.0 182.97 508.44 184.68 ;
   RECT 0.0 184.68 508.44 186.39 ;
   RECT 0.0 186.39 508.44 188.1 ;
   RECT 0.0 188.1 508.44 189.81 ;
   RECT 0.0 189.81 508.44 191.52 ;
   RECT 0.0 191.52 508.44 193.23 ;
   RECT 0.0 193.23 508.44 194.94 ;
   RECT 0.0 194.94 508.44 196.65 ;
   RECT 0.0 196.65 508.44 198.36 ;
   RECT 0.0 198.36 508.44 200.07 ;
   RECT 0.0 200.07 508.44 201.78 ;
   RECT 0.0 201.78 508.44 203.49 ;
   RECT 0.0 203.49 508.44 205.2 ;
   RECT 0.0 205.2 508.44 206.91 ;
   RECT 0.0 206.91 508.44 208.62 ;
   RECT 0.0 208.62 508.44 210.33 ;
   RECT 0.0 210.33 508.44 212.04 ;
   RECT 23.18 212.04 508.44 213.75 ;
   RECT 23.18 213.75 508.44 215.46 ;
   RECT 23.18 215.46 508.44 217.17 ;
   RECT 23.18 217.17 508.44 218.88 ;
   RECT 23.18 218.88 508.44 220.59 ;
   RECT 23.18 220.59 508.44 222.3 ;
   RECT 23.18 222.3 508.44 224.01 ;
   RECT 23.18 224.01 508.44 225.72 ;
   RECT 23.18 225.72 508.44 227.43 ;
   RECT 23.18 227.43 508.44 229.14 ;
   RECT 23.18 229.14 508.44 230.85 ;
   RECT 23.18 230.85 508.44 232.56 ;
   RECT 23.18 232.56 508.44 234.27 ;
   RECT 23.18 234.27 508.44 235.98 ;
   RECT 23.18 235.98 508.44 237.69 ;
   RECT 23.18 237.69 508.44 239.4 ;
   RECT 23.18 239.4 508.44 241.11 ;
   RECT 23.18 241.11 508.44 242.82 ;
   RECT 23.18 242.82 508.44 244.53 ;
   RECT 23.18 244.53 508.44 246.24 ;
   RECT 23.18 246.24 508.44 247.95 ;
   RECT 23.18 247.95 508.44 249.66 ;
   RECT 23.18 249.66 508.44 251.37 ;
   RECT 23.18 251.37 508.44 253.08 ;
   RECT 23.18 253.08 508.44 254.79 ;
   RECT 23.18 254.79 508.44 256.5 ;
   RECT 23.18 256.5 508.44 258.21 ;
   RECT 23.18 258.21 508.44 259.92 ;
   RECT 23.18 259.92 508.44 261.63 ;
   RECT 23.18 261.63 508.44 263.34 ;
   RECT 23.18 263.34 508.44 265.05 ;
   RECT 23.18 265.05 508.44 266.76 ;
   RECT 23.18 266.76 508.44 268.47 ;
   RECT 23.18 268.47 508.44 270.18 ;
   RECT 23.18 270.18 508.44 271.89 ;
   RECT 23.18 271.89 508.44 273.6 ;
   RECT 23.18 273.6 508.44 275.31 ;
   RECT 23.18 275.31 508.44 277.02 ;
   RECT 23.18 277.02 508.44 278.73 ;
   RECT 23.18 278.73 508.44 280.44 ;
   RECT 23.18 280.44 508.44 282.15 ;
   RECT 23.18 282.15 508.44 283.86 ;
   RECT 23.18 283.86 508.44 285.57 ;
   RECT 23.18 285.57 508.44 287.28 ;
   RECT 23.18 287.28 508.44 288.99 ;
   RECT 23.18 288.99 508.44 290.7 ;
   RECT 23.18 290.7 508.44 292.41 ;
   RECT 23.18 292.41 508.44 294.12 ;
   RECT 23.18 294.12 508.44 295.83 ;
   RECT 23.18 295.83 508.44 297.54 ;
   RECT 23.18 297.54 508.44 299.25 ;
   RECT 23.18 299.25 508.44 300.96 ;
   RECT 23.18 300.96 508.44 302.67 ;
   RECT 23.18 302.67 508.44 304.38 ;
   RECT 23.18 304.38 508.44 306.09 ;
   RECT 23.18 306.09 508.44 307.8 ;
   RECT 23.18 307.8 508.44 309.51 ;
   RECT 23.18 309.51 508.44 311.22 ;
   RECT 23.18 311.22 508.44 312.93 ;
   RECT 23.18 312.93 508.44 314.64 ;
   RECT 23.18 314.64 508.44 316.35 ;
   RECT 23.18 316.35 508.44 318.06 ;
   RECT 23.18 318.06 508.44 319.77 ;
   RECT 23.18 319.77 508.44 321.48 ;
   RECT 23.18 321.48 508.44 323.19 ;
   RECT 23.18 323.19 508.44 324.9 ;
   RECT 23.18 324.9 508.44 326.61 ;
   RECT 23.18 326.61 508.44 328.32 ;
   RECT 23.18 328.32 508.44 330.03 ;
   RECT 23.18 330.03 508.44 331.74 ;
   RECT 23.18 331.74 508.44 333.45 ;
   RECT 23.18 333.45 508.44 335.16 ;
   RECT 23.18 335.16 508.44 336.87 ;
   RECT 23.18 336.87 508.44 338.58 ;
   RECT 23.18 338.58 508.44 340.29 ;
   RECT 23.18 340.29 508.44 342.0 ;
   RECT 23.18 342.0 508.44 343.71 ;
   RECT 23.18 343.71 508.44 345.42 ;
   RECT 23.18 345.42 508.44 347.13 ;
   RECT 23.18 347.13 508.44 348.84 ;
   RECT 23.18 348.84 508.44 350.55 ;
   RECT 23.18 350.55 508.44 352.26 ;
   RECT 23.18 352.26 508.44 353.97 ;
   RECT 23.18 353.97 508.44 355.68 ;
   RECT 23.18 355.68 508.44 357.39 ;
   RECT 23.18 357.39 508.44 359.1 ;
   RECT 23.18 359.1 508.44 360.81 ;
   RECT 23.18 360.81 508.44 362.52 ;
   RECT 23.18 362.52 508.44 364.23 ;
   RECT 23.18 364.23 508.44 365.94 ;
   RECT 23.18 365.94 508.44 367.65 ;
   RECT 23.18 367.65 508.44 369.36 ;
   RECT 23.18 369.36 508.44 371.07 ;
   RECT 23.18 371.07 508.44 372.78 ;
   RECT 23.18 372.78 508.44 374.49 ;
   RECT 23.18 374.49 508.44 376.2 ;
   RECT 23.18 376.2 508.44 377.91 ;
   RECT 23.18 377.91 508.44 379.62 ;
   RECT 23.18 379.62 508.44 381.33 ;
   RECT 23.18 381.33 508.44 383.04 ;
   RECT 23.18 383.04 508.44 384.75 ;
   RECT 23.18 384.75 508.44 386.46 ;
   RECT 23.18 386.46 508.44 388.17 ;
   RECT 23.18 388.17 508.44 389.88 ;
   RECT 23.18 389.88 508.44 391.59 ;
   RECT 23.18 391.59 508.44 393.3 ;
   RECT 23.18 393.3 508.44 395.01 ;
   RECT 23.18 395.01 508.44 396.72 ;
   RECT 23.18 396.72 508.44 398.43 ;
   RECT 23.18 398.43 508.44 400.14 ;
   RECT 23.18 400.14 508.44 401.85 ;
   RECT 23.18 401.85 508.44 403.56 ;
   RECT 23.18 403.56 508.44 405.27 ;
   RECT 23.18 405.27 508.44 406.98 ;
   RECT 23.18 406.98 508.44 408.69 ;
   RECT 23.18 408.69 508.44 410.4 ;
  LAYER via2 ;
   RECT 23.18 0.0 508.44 1.71 ;
   RECT 23.18 1.71 508.44 3.42 ;
   RECT 23.18 3.42 508.44 5.13 ;
   RECT 23.18 5.13 508.44 6.84 ;
   RECT 23.18 6.84 508.44 8.55 ;
   RECT 23.18 8.55 508.44 10.26 ;
   RECT 23.18 10.26 508.44 11.97 ;
   RECT 23.18 11.97 508.44 13.68 ;
   RECT 23.18 13.68 508.44 15.39 ;
   RECT 23.18 15.39 508.44 17.1 ;
   RECT 23.18 17.1 508.44 18.81 ;
   RECT 23.18 18.81 508.44 20.52 ;
   RECT 23.18 20.52 508.44 22.23 ;
   RECT 23.18 22.23 508.44 23.94 ;
   RECT 23.18 23.94 508.44 25.65 ;
   RECT 23.18 25.65 508.44 27.36 ;
   RECT 23.18 27.36 508.44 29.07 ;
   RECT 23.18 29.07 508.44 30.78 ;
   RECT 23.18 30.78 508.44 32.49 ;
   RECT 23.18 32.49 508.44 34.2 ;
   RECT 23.18 34.2 508.44 35.91 ;
   RECT 23.18 35.91 508.44 37.62 ;
   RECT 23.18 37.62 508.44 39.33 ;
   RECT 23.18 39.33 508.44 41.04 ;
   RECT 23.18 41.04 508.44 42.75 ;
   RECT 23.18 42.75 508.44 44.46 ;
   RECT 23.18 44.46 508.44 46.17 ;
   RECT 23.18 46.17 508.44 47.88 ;
   RECT 23.18 47.88 508.44 49.59 ;
   RECT 23.18 49.59 508.44 51.3 ;
   RECT 23.18 51.3 508.44 53.01 ;
   RECT 23.18 53.01 508.44 54.72 ;
   RECT 23.18 54.72 508.44 56.43 ;
   RECT 23.18 56.43 508.44 58.14 ;
   RECT 23.18 58.14 508.44 59.85 ;
   RECT 23.18 59.85 508.44 61.56 ;
   RECT 23.18 61.56 508.44 63.27 ;
   RECT 23.18 63.27 508.44 64.98 ;
   RECT 23.18 64.98 508.44 66.69 ;
   RECT 23.18 66.69 508.44 68.4 ;
   RECT 23.18 68.4 508.44 70.11 ;
   RECT 23.18 70.11 508.44 71.82 ;
   RECT 23.18 71.82 508.44 73.53 ;
   RECT 23.18 73.53 508.44 75.24 ;
   RECT 23.18 75.24 508.44 76.95 ;
   RECT 23.18 76.95 508.44 78.66 ;
   RECT 23.18 78.66 508.44 80.37 ;
   RECT 23.18 80.37 508.44 82.08 ;
   RECT 23.18 82.08 508.44 83.79 ;
   RECT 23.18 83.79 508.44 85.5 ;
   RECT 23.18 85.5 508.44 87.21 ;
   RECT 23.18 87.21 508.44 88.92 ;
   RECT 23.18 88.92 508.44 90.63 ;
   RECT 23.18 90.63 508.44 92.34 ;
   RECT 23.18 92.34 508.44 94.05 ;
   RECT 23.18 94.05 508.44 95.76 ;
   RECT 23.18 95.76 508.44 97.47 ;
   RECT 23.18 97.47 508.44 99.18 ;
   RECT 23.18 99.18 508.44 100.89 ;
   RECT 23.18 100.89 508.44 102.6 ;
   RECT 23.18 102.6 508.44 104.31 ;
   RECT 23.18 104.31 508.44 106.02 ;
   RECT 23.18 106.02 508.44 107.73 ;
   RECT 23.18 107.73 508.44 109.44 ;
   RECT 23.18 109.44 508.44 111.15 ;
   RECT 23.18 111.15 508.44 112.86 ;
   RECT 23.18 112.86 508.44 114.57 ;
   RECT 23.18 114.57 508.44 116.28 ;
   RECT 23.18 116.28 508.44 117.99 ;
   RECT 23.18 117.99 508.44 119.7 ;
   RECT 23.18 119.7 508.44 121.41 ;
   RECT 23.18 121.41 508.44 123.12 ;
   RECT 23.18 123.12 508.44 124.83 ;
   RECT 23.18 124.83 508.44 126.54 ;
   RECT 23.18 126.54 508.44 128.25 ;
   RECT 23.18 128.25 508.44 129.96 ;
   RECT 23.18 129.96 508.44 131.67 ;
   RECT 23.18 131.67 508.44 133.38 ;
   RECT 23.18 133.38 508.44 135.09 ;
   RECT 23.18 135.09 508.44 136.8 ;
   RECT 23.18 136.8 508.44 138.51 ;
   RECT 23.18 138.51 508.44 140.22 ;
   RECT 23.18 140.22 508.44 141.93 ;
   RECT 23.18 141.93 508.44 143.64 ;
   RECT 23.18 143.64 508.44 145.35 ;
   RECT 23.18 145.35 508.44 147.06 ;
   RECT 23.18 147.06 508.44 148.77 ;
   RECT 23.18 148.77 508.44 150.48 ;
   RECT 23.18 150.48 508.44 152.19 ;
   RECT 23.18 152.19 508.44 153.9 ;
   RECT 23.18 153.9 508.44 155.61 ;
   RECT 23.18 155.61 508.44 157.32 ;
   RECT 23.18 157.32 508.44 159.03 ;
   RECT 23.18 159.03 508.44 160.74 ;
   RECT 23.18 160.74 508.44 162.45 ;
   RECT 23.18 162.45 508.44 164.16 ;
   RECT 23.18 164.16 508.44 165.87 ;
   RECT 23.18 165.87 508.44 167.58 ;
   RECT 23.18 167.58 508.44 169.29 ;
   RECT 23.18 169.29 508.44 171.0 ;
   RECT 23.18 171.0 508.44 172.71 ;
   RECT 23.18 172.71 508.44 174.42 ;
   RECT 23.18 174.42 508.44 176.13 ;
   RECT 23.18 176.13 508.44 177.84 ;
   RECT 23.18 177.84 508.44 179.55 ;
   RECT 23.18 179.55 508.44 181.26 ;
   RECT 23.18 181.26 508.44 182.97 ;
   RECT 0.0 182.97 508.44 184.68 ;
   RECT 0.0 184.68 508.44 186.39 ;
   RECT 0.0 186.39 508.44 188.1 ;
   RECT 0.0 188.1 508.44 189.81 ;
   RECT 0.0 189.81 508.44 191.52 ;
   RECT 0.0 191.52 508.44 193.23 ;
   RECT 0.0 193.23 508.44 194.94 ;
   RECT 0.0 194.94 508.44 196.65 ;
   RECT 0.0 196.65 508.44 198.36 ;
   RECT 0.0 198.36 508.44 200.07 ;
   RECT 0.0 200.07 508.44 201.78 ;
   RECT 0.0 201.78 508.44 203.49 ;
   RECT 0.0 203.49 508.44 205.2 ;
   RECT 0.0 205.2 508.44 206.91 ;
   RECT 0.0 206.91 508.44 208.62 ;
   RECT 0.0 208.62 508.44 210.33 ;
   RECT 0.0 210.33 508.44 212.04 ;
   RECT 23.18 212.04 508.44 213.75 ;
   RECT 23.18 213.75 508.44 215.46 ;
   RECT 23.18 215.46 508.44 217.17 ;
   RECT 23.18 217.17 508.44 218.88 ;
   RECT 23.18 218.88 508.44 220.59 ;
   RECT 23.18 220.59 508.44 222.3 ;
   RECT 23.18 222.3 508.44 224.01 ;
   RECT 23.18 224.01 508.44 225.72 ;
   RECT 23.18 225.72 508.44 227.43 ;
   RECT 23.18 227.43 508.44 229.14 ;
   RECT 23.18 229.14 508.44 230.85 ;
   RECT 23.18 230.85 508.44 232.56 ;
   RECT 23.18 232.56 508.44 234.27 ;
   RECT 23.18 234.27 508.44 235.98 ;
   RECT 23.18 235.98 508.44 237.69 ;
   RECT 23.18 237.69 508.44 239.4 ;
   RECT 23.18 239.4 508.44 241.11 ;
   RECT 23.18 241.11 508.44 242.82 ;
   RECT 23.18 242.82 508.44 244.53 ;
   RECT 23.18 244.53 508.44 246.24 ;
   RECT 23.18 246.24 508.44 247.95 ;
   RECT 23.18 247.95 508.44 249.66 ;
   RECT 23.18 249.66 508.44 251.37 ;
   RECT 23.18 251.37 508.44 253.08 ;
   RECT 23.18 253.08 508.44 254.79 ;
   RECT 23.18 254.79 508.44 256.5 ;
   RECT 23.18 256.5 508.44 258.21 ;
   RECT 23.18 258.21 508.44 259.92 ;
   RECT 23.18 259.92 508.44 261.63 ;
   RECT 23.18 261.63 508.44 263.34 ;
   RECT 23.18 263.34 508.44 265.05 ;
   RECT 23.18 265.05 508.44 266.76 ;
   RECT 23.18 266.76 508.44 268.47 ;
   RECT 23.18 268.47 508.44 270.18 ;
   RECT 23.18 270.18 508.44 271.89 ;
   RECT 23.18 271.89 508.44 273.6 ;
   RECT 23.18 273.6 508.44 275.31 ;
   RECT 23.18 275.31 508.44 277.02 ;
   RECT 23.18 277.02 508.44 278.73 ;
   RECT 23.18 278.73 508.44 280.44 ;
   RECT 23.18 280.44 508.44 282.15 ;
   RECT 23.18 282.15 508.44 283.86 ;
   RECT 23.18 283.86 508.44 285.57 ;
   RECT 23.18 285.57 508.44 287.28 ;
   RECT 23.18 287.28 508.44 288.99 ;
   RECT 23.18 288.99 508.44 290.7 ;
   RECT 23.18 290.7 508.44 292.41 ;
   RECT 23.18 292.41 508.44 294.12 ;
   RECT 23.18 294.12 508.44 295.83 ;
   RECT 23.18 295.83 508.44 297.54 ;
   RECT 23.18 297.54 508.44 299.25 ;
   RECT 23.18 299.25 508.44 300.96 ;
   RECT 23.18 300.96 508.44 302.67 ;
   RECT 23.18 302.67 508.44 304.38 ;
   RECT 23.18 304.38 508.44 306.09 ;
   RECT 23.18 306.09 508.44 307.8 ;
   RECT 23.18 307.8 508.44 309.51 ;
   RECT 23.18 309.51 508.44 311.22 ;
   RECT 23.18 311.22 508.44 312.93 ;
   RECT 23.18 312.93 508.44 314.64 ;
   RECT 23.18 314.64 508.44 316.35 ;
   RECT 23.18 316.35 508.44 318.06 ;
   RECT 23.18 318.06 508.44 319.77 ;
   RECT 23.18 319.77 508.44 321.48 ;
   RECT 23.18 321.48 508.44 323.19 ;
   RECT 23.18 323.19 508.44 324.9 ;
   RECT 23.18 324.9 508.44 326.61 ;
   RECT 23.18 326.61 508.44 328.32 ;
   RECT 23.18 328.32 508.44 330.03 ;
   RECT 23.18 330.03 508.44 331.74 ;
   RECT 23.18 331.74 508.44 333.45 ;
   RECT 23.18 333.45 508.44 335.16 ;
   RECT 23.18 335.16 508.44 336.87 ;
   RECT 23.18 336.87 508.44 338.58 ;
   RECT 23.18 338.58 508.44 340.29 ;
   RECT 23.18 340.29 508.44 342.0 ;
   RECT 23.18 342.0 508.44 343.71 ;
   RECT 23.18 343.71 508.44 345.42 ;
   RECT 23.18 345.42 508.44 347.13 ;
   RECT 23.18 347.13 508.44 348.84 ;
   RECT 23.18 348.84 508.44 350.55 ;
   RECT 23.18 350.55 508.44 352.26 ;
   RECT 23.18 352.26 508.44 353.97 ;
   RECT 23.18 353.97 508.44 355.68 ;
   RECT 23.18 355.68 508.44 357.39 ;
   RECT 23.18 357.39 508.44 359.1 ;
   RECT 23.18 359.1 508.44 360.81 ;
   RECT 23.18 360.81 508.44 362.52 ;
   RECT 23.18 362.52 508.44 364.23 ;
   RECT 23.18 364.23 508.44 365.94 ;
   RECT 23.18 365.94 508.44 367.65 ;
   RECT 23.18 367.65 508.44 369.36 ;
   RECT 23.18 369.36 508.44 371.07 ;
   RECT 23.18 371.07 508.44 372.78 ;
   RECT 23.18 372.78 508.44 374.49 ;
   RECT 23.18 374.49 508.44 376.2 ;
   RECT 23.18 376.2 508.44 377.91 ;
   RECT 23.18 377.91 508.44 379.62 ;
   RECT 23.18 379.62 508.44 381.33 ;
   RECT 23.18 381.33 508.44 383.04 ;
   RECT 23.18 383.04 508.44 384.75 ;
   RECT 23.18 384.75 508.44 386.46 ;
   RECT 23.18 386.46 508.44 388.17 ;
   RECT 23.18 388.17 508.44 389.88 ;
   RECT 23.18 389.88 508.44 391.59 ;
   RECT 23.18 391.59 508.44 393.3 ;
   RECT 23.18 393.3 508.44 395.01 ;
   RECT 23.18 395.01 508.44 396.72 ;
   RECT 23.18 396.72 508.44 398.43 ;
   RECT 23.18 398.43 508.44 400.14 ;
   RECT 23.18 400.14 508.44 401.85 ;
   RECT 23.18 401.85 508.44 403.56 ;
   RECT 23.18 403.56 508.44 405.27 ;
   RECT 23.18 405.27 508.44 406.98 ;
   RECT 23.18 406.98 508.44 408.69 ;
   RECT 23.18 408.69 508.44 410.4 ;
  LAYER metal3 ;
   RECT 23.18 0.0 508.44 1.71 ;
   RECT 23.18 1.71 508.44 3.42 ;
   RECT 23.18 3.42 508.44 5.13 ;
   RECT 23.18 5.13 508.44 6.84 ;
   RECT 23.18 6.84 508.44 8.55 ;
   RECT 23.18 8.55 508.44 10.26 ;
   RECT 23.18 10.26 508.44 11.97 ;
   RECT 23.18 11.97 508.44 13.68 ;
   RECT 23.18 13.68 508.44 15.39 ;
   RECT 23.18 15.39 508.44 17.1 ;
   RECT 23.18 17.1 508.44 18.81 ;
   RECT 23.18 18.81 508.44 20.52 ;
   RECT 23.18 20.52 508.44 22.23 ;
   RECT 23.18 22.23 508.44 23.94 ;
   RECT 23.18 23.94 508.44 25.65 ;
   RECT 23.18 25.65 508.44 27.36 ;
   RECT 23.18 27.36 508.44 29.07 ;
   RECT 23.18 29.07 508.44 30.78 ;
   RECT 23.18 30.78 508.44 32.49 ;
   RECT 23.18 32.49 508.44 34.2 ;
   RECT 23.18 34.2 508.44 35.91 ;
   RECT 23.18 35.91 508.44 37.62 ;
   RECT 23.18 37.62 508.44 39.33 ;
   RECT 23.18 39.33 508.44 41.04 ;
   RECT 23.18 41.04 508.44 42.75 ;
   RECT 23.18 42.75 508.44 44.46 ;
   RECT 23.18 44.46 508.44 46.17 ;
   RECT 23.18 46.17 508.44 47.88 ;
   RECT 23.18 47.88 508.44 49.59 ;
   RECT 23.18 49.59 508.44 51.3 ;
   RECT 23.18 51.3 508.44 53.01 ;
   RECT 23.18 53.01 508.44 54.72 ;
   RECT 23.18 54.72 508.44 56.43 ;
   RECT 23.18 56.43 508.44 58.14 ;
   RECT 23.18 58.14 508.44 59.85 ;
   RECT 23.18 59.85 508.44 61.56 ;
   RECT 23.18 61.56 508.44 63.27 ;
   RECT 23.18 63.27 508.44 64.98 ;
   RECT 23.18 64.98 508.44 66.69 ;
   RECT 23.18 66.69 508.44 68.4 ;
   RECT 23.18 68.4 508.44 70.11 ;
   RECT 23.18 70.11 508.44 71.82 ;
   RECT 23.18 71.82 508.44 73.53 ;
   RECT 23.18 73.53 508.44 75.24 ;
   RECT 23.18 75.24 508.44 76.95 ;
   RECT 23.18 76.95 508.44 78.66 ;
   RECT 23.18 78.66 508.44 80.37 ;
   RECT 23.18 80.37 508.44 82.08 ;
   RECT 23.18 82.08 508.44 83.79 ;
   RECT 23.18 83.79 508.44 85.5 ;
   RECT 23.18 85.5 508.44 87.21 ;
   RECT 23.18 87.21 508.44 88.92 ;
   RECT 23.18 88.92 508.44 90.63 ;
   RECT 23.18 90.63 508.44 92.34 ;
   RECT 23.18 92.34 508.44 94.05 ;
   RECT 23.18 94.05 508.44 95.76 ;
   RECT 23.18 95.76 508.44 97.47 ;
   RECT 23.18 97.47 508.44 99.18 ;
   RECT 23.18 99.18 508.44 100.89 ;
   RECT 23.18 100.89 508.44 102.6 ;
   RECT 23.18 102.6 508.44 104.31 ;
   RECT 23.18 104.31 508.44 106.02 ;
   RECT 23.18 106.02 508.44 107.73 ;
   RECT 23.18 107.73 508.44 109.44 ;
   RECT 23.18 109.44 508.44 111.15 ;
   RECT 23.18 111.15 508.44 112.86 ;
   RECT 23.18 112.86 508.44 114.57 ;
   RECT 23.18 114.57 508.44 116.28 ;
   RECT 23.18 116.28 508.44 117.99 ;
   RECT 23.18 117.99 508.44 119.7 ;
   RECT 23.18 119.7 508.44 121.41 ;
   RECT 23.18 121.41 508.44 123.12 ;
   RECT 23.18 123.12 508.44 124.83 ;
   RECT 23.18 124.83 508.44 126.54 ;
   RECT 23.18 126.54 508.44 128.25 ;
   RECT 23.18 128.25 508.44 129.96 ;
   RECT 23.18 129.96 508.44 131.67 ;
   RECT 23.18 131.67 508.44 133.38 ;
   RECT 23.18 133.38 508.44 135.09 ;
   RECT 23.18 135.09 508.44 136.8 ;
   RECT 23.18 136.8 508.44 138.51 ;
   RECT 23.18 138.51 508.44 140.22 ;
   RECT 23.18 140.22 508.44 141.93 ;
   RECT 23.18 141.93 508.44 143.64 ;
   RECT 23.18 143.64 508.44 145.35 ;
   RECT 23.18 145.35 508.44 147.06 ;
   RECT 23.18 147.06 508.44 148.77 ;
   RECT 23.18 148.77 508.44 150.48 ;
   RECT 23.18 150.48 508.44 152.19 ;
   RECT 23.18 152.19 508.44 153.9 ;
   RECT 23.18 153.9 508.44 155.61 ;
   RECT 23.18 155.61 508.44 157.32 ;
   RECT 23.18 157.32 508.44 159.03 ;
   RECT 23.18 159.03 508.44 160.74 ;
   RECT 23.18 160.74 508.44 162.45 ;
   RECT 23.18 162.45 508.44 164.16 ;
   RECT 23.18 164.16 508.44 165.87 ;
   RECT 23.18 165.87 508.44 167.58 ;
   RECT 23.18 167.58 508.44 169.29 ;
   RECT 23.18 169.29 508.44 171.0 ;
   RECT 23.18 171.0 508.44 172.71 ;
   RECT 23.18 172.71 508.44 174.42 ;
   RECT 23.18 174.42 508.44 176.13 ;
   RECT 23.18 176.13 508.44 177.84 ;
   RECT 23.18 177.84 508.44 179.55 ;
   RECT 23.18 179.55 508.44 181.26 ;
   RECT 23.18 181.26 508.44 182.97 ;
   RECT 0.0 182.97 508.44 184.68 ;
   RECT 0.0 184.68 508.44 186.39 ;
   RECT 0.0 186.39 508.44 188.1 ;
   RECT 0.0 188.1 508.44 189.81 ;
   RECT 0.0 189.81 508.44 191.52 ;
   RECT 0.0 191.52 508.44 193.23 ;
   RECT 0.0 193.23 508.44 194.94 ;
   RECT 0.0 194.94 508.44 196.65 ;
   RECT 0.0 196.65 508.44 198.36 ;
   RECT 0.0 198.36 508.44 200.07 ;
   RECT 0.0 200.07 508.44 201.78 ;
   RECT 0.0 201.78 508.44 203.49 ;
   RECT 0.0 203.49 508.44 205.2 ;
   RECT 0.0 205.2 508.44 206.91 ;
   RECT 0.0 206.91 508.44 208.62 ;
   RECT 0.0 208.62 508.44 210.33 ;
   RECT 0.0 210.33 508.44 212.04 ;
   RECT 23.18 212.04 508.44 213.75 ;
   RECT 23.18 213.75 508.44 215.46 ;
   RECT 23.18 215.46 508.44 217.17 ;
   RECT 23.18 217.17 508.44 218.88 ;
   RECT 23.18 218.88 508.44 220.59 ;
   RECT 23.18 220.59 508.44 222.3 ;
   RECT 23.18 222.3 508.44 224.01 ;
   RECT 23.18 224.01 508.44 225.72 ;
   RECT 23.18 225.72 508.44 227.43 ;
   RECT 23.18 227.43 508.44 229.14 ;
   RECT 23.18 229.14 508.44 230.85 ;
   RECT 23.18 230.85 508.44 232.56 ;
   RECT 23.18 232.56 508.44 234.27 ;
   RECT 23.18 234.27 508.44 235.98 ;
   RECT 23.18 235.98 508.44 237.69 ;
   RECT 23.18 237.69 508.44 239.4 ;
   RECT 23.18 239.4 508.44 241.11 ;
   RECT 23.18 241.11 508.44 242.82 ;
   RECT 23.18 242.82 508.44 244.53 ;
   RECT 23.18 244.53 508.44 246.24 ;
   RECT 23.18 246.24 508.44 247.95 ;
   RECT 23.18 247.95 508.44 249.66 ;
   RECT 23.18 249.66 508.44 251.37 ;
   RECT 23.18 251.37 508.44 253.08 ;
   RECT 23.18 253.08 508.44 254.79 ;
   RECT 23.18 254.79 508.44 256.5 ;
   RECT 23.18 256.5 508.44 258.21 ;
   RECT 23.18 258.21 508.44 259.92 ;
   RECT 23.18 259.92 508.44 261.63 ;
   RECT 23.18 261.63 508.44 263.34 ;
   RECT 23.18 263.34 508.44 265.05 ;
   RECT 23.18 265.05 508.44 266.76 ;
   RECT 23.18 266.76 508.44 268.47 ;
   RECT 23.18 268.47 508.44 270.18 ;
   RECT 23.18 270.18 508.44 271.89 ;
   RECT 23.18 271.89 508.44 273.6 ;
   RECT 23.18 273.6 508.44 275.31 ;
   RECT 23.18 275.31 508.44 277.02 ;
   RECT 23.18 277.02 508.44 278.73 ;
   RECT 23.18 278.73 508.44 280.44 ;
   RECT 23.18 280.44 508.44 282.15 ;
   RECT 23.18 282.15 508.44 283.86 ;
   RECT 23.18 283.86 508.44 285.57 ;
   RECT 23.18 285.57 508.44 287.28 ;
   RECT 23.18 287.28 508.44 288.99 ;
   RECT 23.18 288.99 508.44 290.7 ;
   RECT 23.18 290.7 508.44 292.41 ;
   RECT 23.18 292.41 508.44 294.12 ;
   RECT 23.18 294.12 508.44 295.83 ;
   RECT 23.18 295.83 508.44 297.54 ;
   RECT 23.18 297.54 508.44 299.25 ;
   RECT 23.18 299.25 508.44 300.96 ;
   RECT 23.18 300.96 508.44 302.67 ;
   RECT 23.18 302.67 508.44 304.38 ;
   RECT 23.18 304.38 508.44 306.09 ;
   RECT 23.18 306.09 508.44 307.8 ;
   RECT 23.18 307.8 508.44 309.51 ;
   RECT 23.18 309.51 508.44 311.22 ;
   RECT 23.18 311.22 508.44 312.93 ;
   RECT 23.18 312.93 508.44 314.64 ;
   RECT 23.18 314.64 508.44 316.35 ;
   RECT 23.18 316.35 508.44 318.06 ;
   RECT 23.18 318.06 508.44 319.77 ;
   RECT 23.18 319.77 508.44 321.48 ;
   RECT 23.18 321.48 508.44 323.19 ;
   RECT 23.18 323.19 508.44 324.9 ;
   RECT 23.18 324.9 508.44 326.61 ;
   RECT 23.18 326.61 508.44 328.32 ;
   RECT 23.18 328.32 508.44 330.03 ;
   RECT 23.18 330.03 508.44 331.74 ;
   RECT 23.18 331.74 508.44 333.45 ;
   RECT 23.18 333.45 508.44 335.16 ;
   RECT 23.18 335.16 508.44 336.87 ;
   RECT 23.18 336.87 508.44 338.58 ;
   RECT 23.18 338.58 508.44 340.29 ;
   RECT 23.18 340.29 508.44 342.0 ;
   RECT 23.18 342.0 508.44 343.71 ;
   RECT 23.18 343.71 508.44 345.42 ;
   RECT 23.18 345.42 508.44 347.13 ;
   RECT 23.18 347.13 508.44 348.84 ;
   RECT 23.18 348.84 508.44 350.55 ;
   RECT 23.18 350.55 508.44 352.26 ;
   RECT 23.18 352.26 508.44 353.97 ;
   RECT 23.18 353.97 508.44 355.68 ;
   RECT 23.18 355.68 508.44 357.39 ;
   RECT 23.18 357.39 508.44 359.1 ;
   RECT 23.18 359.1 508.44 360.81 ;
   RECT 23.18 360.81 508.44 362.52 ;
   RECT 23.18 362.52 508.44 364.23 ;
   RECT 23.18 364.23 508.44 365.94 ;
   RECT 23.18 365.94 508.44 367.65 ;
   RECT 23.18 367.65 508.44 369.36 ;
   RECT 23.18 369.36 508.44 371.07 ;
   RECT 23.18 371.07 508.44 372.78 ;
   RECT 23.18 372.78 508.44 374.49 ;
   RECT 23.18 374.49 508.44 376.2 ;
   RECT 23.18 376.2 508.44 377.91 ;
   RECT 23.18 377.91 508.44 379.62 ;
   RECT 23.18 379.62 508.44 381.33 ;
   RECT 23.18 381.33 508.44 383.04 ;
   RECT 23.18 383.04 508.44 384.75 ;
   RECT 23.18 384.75 508.44 386.46 ;
   RECT 23.18 386.46 508.44 388.17 ;
   RECT 23.18 388.17 508.44 389.88 ;
   RECT 23.18 389.88 508.44 391.59 ;
   RECT 23.18 391.59 508.44 393.3 ;
   RECT 23.18 393.3 508.44 395.01 ;
   RECT 23.18 395.01 508.44 396.72 ;
   RECT 23.18 396.72 508.44 398.43 ;
   RECT 23.18 398.43 508.44 400.14 ;
   RECT 23.18 400.14 508.44 401.85 ;
   RECT 23.18 401.85 508.44 403.56 ;
   RECT 23.18 403.56 508.44 405.27 ;
   RECT 23.18 405.27 508.44 406.98 ;
   RECT 23.18 406.98 508.44 408.69 ;
   RECT 23.18 408.69 508.44 410.4 ;
  LAYER via3 ;
   RECT 23.18 0.0 508.44 1.71 ;
   RECT 23.18 1.71 508.44 3.42 ;
   RECT 23.18 3.42 508.44 5.13 ;
   RECT 23.18 5.13 508.44 6.84 ;
   RECT 23.18 6.84 508.44 8.55 ;
   RECT 23.18 8.55 508.44 10.26 ;
   RECT 23.18 10.26 508.44 11.97 ;
   RECT 23.18 11.97 508.44 13.68 ;
   RECT 23.18 13.68 508.44 15.39 ;
   RECT 23.18 15.39 508.44 17.1 ;
   RECT 23.18 17.1 508.44 18.81 ;
   RECT 23.18 18.81 508.44 20.52 ;
   RECT 23.18 20.52 508.44 22.23 ;
   RECT 23.18 22.23 508.44 23.94 ;
   RECT 23.18 23.94 508.44 25.65 ;
   RECT 23.18 25.65 508.44 27.36 ;
   RECT 23.18 27.36 508.44 29.07 ;
   RECT 23.18 29.07 508.44 30.78 ;
   RECT 23.18 30.78 508.44 32.49 ;
   RECT 23.18 32.49 508.44 34.2 ;
   RECT 23.18 34.2 508.44 35.91 ;
   RECT 23.18 35.91 508.44 37.62 ;
   RECT 23.18 37.62 508.44 39.33 ;
   RECT 23.18 39.33 508.44 41.04 ;
   RECT 23.18 41.04 508.44 42.75 ;
   RECT 23.18 42.75 508.44 44.46 ;
   RECT 23.18 44.46 508.44 46.17 ;
   RECT 23.18 46.17 508.44 47.88 ;
   RECT 23.18 47.88 508.44 49.59 ;
   RECT 23.18 49.59 508.44 51.3 ;
   RECT 23.18 51.3 508.44 53.01 ;
   RECT 23.18 53.01 508.44 54.72 ;
   RECT 23.18 54.72 508.44 56.43 ;
   RECT 23.18 56.43 508.44 58.14 ;
   RECT 23.18 58.14 508.44 59.85 ;
   RECT 23.18 59.85 508.44 61.56 ;
   RECT 23.18 61.56 508.44 63.27 ;
   RECT 23.18 63.27 508.44 64.98 ;
   RECT 23.18 64.98 508.44 66.69 ;
   RECT 23.18 66.69 508.44 68.4 ;
   RECT 23.18 68.4 508.44 70.11 ;
   RECT 23.18 70.11 508.44 71.82 ;
   RECT 23.18 71.82 508.44 73.53 ;
   RECT 23.18 73.53 508.44 75.24 ;
   RECT 23.18 75.24 508.44 76.95 ;
   RECT 23.18 76.95 508.44 78.66 ;
   RECT 23.18 78.66 508.44 80.37 ;
   RECT 23.18 80.37 508.44 82.08 ;
   RECT 23.18 82.08 508.44 83.79 ;
   RECT 23.18 83.79 508.44 85.5 ;
   RECT 23.18 85.5 508.44 87.21 ;
   RECT 23.18 87.21 508.44 88.92 ;
   RECT 23.18 88.92 508.44 90.63 ;
   RECT 23.18 90.63 508.44 92.34 ;
   RECT 23.18 92.34 508.44 94.05 ;
   RECT 23.18 94.05 508.44 95.76 ;
   RECT 23.18 95.76 508.44 97.47 ;
   RECT 23.18 97.47 508.44 99.18 ;
   RECT 23.18 99.18 508.44 100.89 ;
   RECT 23.18 100.89 508.44 102.6 ;
   RECT 23.18 102.6 508.44 104.31 ;
   RECT 23.18 104.31 508.44 106.02 ;
   RECT 23.18 106.02 508.44 107.73 ;
   RECT 23.18 107.73 508.44 109.44 ;
   RECT 23.18 109.44 508.44 111.15 ;
   RECT 23.18 111.15 508.44 112.86 ;
   RECT 23.18 112.86 508.44 114.57 ;
   RECT 23.18 114.57 508.44 116.28 ;
   RECT 23.18 116.28 508.44 117.99 ;
   RECT 23.18 117.99 508.44 119.7 ;
   RECT 23.18 119.7 508.44 121.41 ;
   RECT 23.18 121.41 508.44 123.12 ;
   RECT 23.18 123.12 508.44 124.83 ;
   RECT 23.18 124.83 508.44 126.54 ;
   RECT 23.18 126.54 508.44 128.25 ;
   RECT 23.18 128.25 508.44 129.96 ;
   RECT 23.18 129.96 508.44 131.67 ;
   RECT 23.18 131.67 508.44 133.38 ;
   RECT 23.18 133.38 508.44 135.09 ;
   RECT 23.18 135.09 508.44 136.8 ;
   RECT 23.18 136.8 508.44 138.51 ;
   RECT 23.18 138.51 508.44 140.22 ;
   RECT 23.18 140.22 508.44 141.93 ;
   RECT 23.18 141.93 508.44 143.64 ;
   RECT 23.18 143.64 508.44 145.35 ;
   RECT 23.18 145.35 508.44 147.06 ;
   RECT 23.18 147.06 508.44 148.77 ;
   RECT 23.18 148.77 508.44 150.48 ;
   RECT 23.18 150.48 508.44 152.19 ;
   RECT 23.18 152.19 508.44 153.9 ;
   RECT 23.18 153.9 508.44 155.61 ;
   RECT 23.18 155.61 508.44 157.32 ;
   RECT 23.18 157.32 508.44 159.03 ;
   RECT 23.18 159.03 508.44 160.74 ;
   RECT 23.18 160.74 508.44 162.45 ;
   RECT 23.18 162.45 508.44 164.16 ;
   RECT 23.18 164.16 508.44 165.87 ;
   RECT 23.18 165.87 508.44 167.58 ;
   RECT 23.18 167.58 508.44 169.29 ;
   RECT 23.18 169.29 508.44 171.0 ;
   RECT 23.18 171.0 508.44 172.71 ;
   RECT 23.18 172.71 508.44 174.42 ;
   RECT 23.18 174.42 508.44 176.13 ;
   RECT 23.18 176.13 508.44 177.84 ;
   RECT 23.18 177.84 508.44 179.55 ;
   RECT 23.18 179.55 508.44 181.26 ;
   RECT 23.18 181.26 508.44 182.97 ;
   RECT 0.0 182.97 508.44 184.68 ;
   RECT 0.0 184.68 508.44 186.39 ;
   RECT 0.0 186.39 508.44 188.1 ;
   RECT 0.0 188.1 508.44 189.81 ;
   RECT 0.0 189.81 508.44 191.52 ;
   RECT 0.0 191.52 508.44 193.23 ;
   RECT 0.0 193.23 508.44 194.94 ;
   RECT 0.0 194.94 508.44 196.65 ;
   RECT 0.0 196.65 508.44 198.36 ;
   RECT 0.0 198.36 508.44 200.07 ;
   RECT 0.0 200.07 508.44 201.78 ;
   RECT 0.0 201.78 508.44 203.49 ;
   RECT 0.0 203.49 508.44 205.2 ;
   RECT 0.0 205.2 508.44 206.91 ;
   RECT 0.0 206.91 508.44 208.62 ;
   RECT 0.0 208.62 508.44 210.33 ;
   RECT 0.0 210.33 508.44 212.04 ;
   RECT 23.18 212.04 508.44 213.75 ;
   RECT 23.18 213.75 508.44 215.46 ;
   RECT 23.18 215.46 508.44 217.17 ;
   RECT 23.18 217.17 508.44 218.88 ;
   RECT 23.18 218.88 508.44 220.59 ;
   RECT 23.18 220.59 508.44 222.3 ;
   RECT 23.18 222.3 508.44 224.01 ;
   RECT 23.18 224.01 508.44 225.72 ;
   RECT 23.18 225.72 508.44 227.43 ;
   RECT 23.18 227.43 508.44 229.14 ;
   RECT 23.18 229.14 508.44 230.85 ;
   RECT 23.18 230.85 508.44 232.56 ;
   RECT 23.18 232.56 508.44 234.27 ;
   RECT 23.18 234.27 508.44 235.98 ;
   RECT 23.18 235.98 508.44 237.69 ;
   RECT 23.18 237.69 508.44 239.4 ;
   RECT 23.18 239.4 508.44 241.11 ;
   RECT 23.18 241.11 508.44 242.82 ;
   RECT 23.18 242.82 508.44 244.53 ;
   RECT 23.18 244.53 508.44 246.24 ;
   RECT 23.18 246.24 508.44 247.95 ;
   RECT 23.18 247.95 508.44 249.66 ;
   RECT 23.18 249.66 508.44 251.37 ;
   RECT 23.18 251.37 508.44 253.08 ;
   RECT 23.18 253.08 508.44 254.79 ;
   RECT 23.18 254.79 508.44 256.5 ;
   RECT 23.18 256.5 508.44 258.21 ;
   RECT 23.18 258.21 508.44 259.92 ;
   RECT 23.18 259.92 508.44 261.63 ;
   RECT 23.18 261.63 508.44 263.34 ;
   RECT 23.18 263.34 508.44 265.05 ;
   RECT 23.18 265.05 508.44 266.76 ;
   RECT 23.18 266.76 508.44 268.47 ;
   RECT 23.18 268.47 508.44 270.18 ;
   RECT 23.18 270.18 508.44 271.89 ;
   RECT 23.18 271.89 508.44 273.6 ;
   RECT 23.18 273.6 508.44 275.31 ;
   RECT 23.18 275.31 508.44 277.02 ;
   RECT 23.18 277.02 508.44 278.73 ;
   RECT 23.18 278.73 508.44 280.44 ;
   RECT 23.18 280.44 508.44 282.15 ;
   RECT 23.18 282.15 508.44 283.86 ;
   RECT 23.18 283.86 508.44 285.57 ;
   RECT 23.18 285.57 508.44 287.28 ;
   RECT 23.18 287.28 508.44 288.99 ;
   RECT 23.18 288.99 508.44 290.7 ;
   RECT 23.18 290.7 508.44 292.41 ;
   RECT 23.18 292.41 508.44 294.12 ;
   RECT 23.18 294.12 508.44 295.83 ;
   RECT 23.18 295.83 508.44 297.54 ;
   RECT 23.18 297.54 508.44 299.25 ;
   RECT 23.18 299.25 508.44 300.96 ;
   RECT 23.18 300.96 508.44 302.67 ;
   RECT 23.18 302.67 508.44 304.38 ;
   RECT 23.18 304.38 508.44 306.09 ;
   RECT 23.18 306.09 508.44 307.8 ;
   RECT 23.18 307.8 508.44 309.51 ;
   RECT 23.18 309.51 508.44 311.22 ;
   RECT 23.18 311.22 508.44 312.93 ;
   RECT 23.18 312.93 508.44 314.64 ;
   RECT 23.18 314.64 508.44 316.35 ;
   RECT 23.18 316.35 508.44 318.06 ;
   RECT 23.18 318.06 508.44 319.77 ;
   RECT 23.18 319.77 508.44 321.48 ;
   RECT 23.18 321.48 508.44 323.19 ;
   RECT 23.18 323.19 508.44 324.9 ;
   RECT 23.18 324.9 508.44 326.61 ;
   RECT 23.18 326.61 508.44 328.32 ;
   RECT 23.18 328.32 508.44 330.03 ;
   RECT 23.18 330.03 508.44 331.74 ;
   RECT 23.18 331.74 508.44 333.45 ;
   RECT 23.18 333.45 508.44 335.16 ;
   RECT 23.18 335.16 508.44 336.87 ;
   RECT 23.18 336.87 508.44 338.58 ;
   RECT 23.18 338.58 508.44 340.29 ;
   RECT 23.18 340.29 508.44 342.0 ;
   RECT 23.18 342.0 508.44 343.71 ;
   RECT 23.18 343.71 508.44 345.42 ;
   RECT 23.18 345.42 508.44 347.13 ;
   RECT 23.18 347.13 508.44 348.84 ;
   RECT 23.18 348.84 508.44 350.55 ;
   RECT 23.18 350.55 508.44 352.26 ;
   RECT 23.18 352.26 508.44 353.97 ;
   RECT 23.18 353.97 508.44 355.68 ;
   RECT 23.18 355.68 508.44 357.39 ;
   RECT 23.18 357.39 508.44 359.1 ;
   RECT 23.18 359.1 508.44 360.81 ;
   RECT 23.18 360.81 508.44 362.52 ;
   RECT 23.18 362.52 508.44 364.23 ;
   RECT 23.18 364.23 508.44 365.94 ;
   RECT 23.18 365.94 508.44 367.65 ;
   RECT 23.18 367.65 508.44 369.36 ;
   RECT 23.18 369.36 508.44 371.07 ;
   RECT 23.18 371.07 508.44 372.78 ;
   RECT 23.18 372.78 508.44 374.49 ;
   RECT 23.18 374.49 508.44 376.2 ;
   RECT 23.18 376.2 508.44 377.91 ;
   RECT 23.18 377.91 508.44 379.62 ;
   RECT 23.18 379.62 508.44 381.33 ;
   RECT 23.18 381.33 508.44 383.04 ;
   RECT 23.18 383.04 508.44 384.75 ;
   RECT 23.18 384.75 508.44 386.46 ;
   RECT 23.18 386.46 508.44 388.17 ;
   RECT 23.18 388.17 508.44 389.88 ;
   RECT 23.18 389.88 508.44 391.59 ;
   RECT 23.18 391.59 508.44 393.3 ;
   RECT 23.18 393.3 508.44 395.01 ;
   RECT 23.18 395.01 508.44 396.72 ;
   RECT 23.18 396.72 508.44 398.43 ;
   RECT 23.18 398.43 508.44 400.14 ;
   RECT 23.18 400.14 508.44 401.85 ;
   RECT 23.18 401.85 508.44 403.56 ;
   RECT 23.18 403.56 508.44 405.27 ;
   RECT 23.18 405.27 508.44 406.98 ;
   RECT 23.18 406.98 508.44 408.69 ;
   RECT 23.18 408.69 508.44 410.4 ;
  LAYER metal4 ;
   RECT 23.18 0.0 508.44 1.71 ;
   RECT 23.18 1.71 508.44 3.42 ;
   RECT 23.18 3.42 508.44 5.13 ;
   RECT 23.18 5.13 508.44 6.84 ;
   RECT 23.18 6.84 508.44 8.55 ;
   RECT 23.18 8.55 508.44 10.26 ;
   RECT 23.18 10.26 508.44 11.97 ;
   RECT 23.18 11.97 508.44 13.68 ;
   RECT 23.18 13.68 508.44 15.39 ;
   RECT 23.18 15.39 508.44 17.1 ;
   RECT 23.18 17.1 508.44 18.81 ;
   RECT 23.18 18.81 508.44 20.52 ;
   RECT 23.18 20.52 508.44 22.23 ;
   RECT 23.18 22.23 508.44 23.94 ;
   RECT 23.18 23.94 508.44 25.65 ;
   RECT 23.18 25.65 508.44 27.36 ;
   RECT 23.18 27.36 508.44 29.07 ;
   RECT 23.18 29.07 508.44 30.78 ;
   RECT 23.18 30.78 508.44 32.49 ;
   RECT 23.18 32.49 508.44 34.2 ;
   RECT 23.18 34.2 508.44 35.91 ;
   RECT 23.18 35.91 508.44 37.62 ;
   RECT 23.18 37.62 508.44 39.33 ;
   RECT 23.18 39.33 508.44 41.04 ;
   RECT 23.18 41.04 508.44 42.75 ;
   RECT 23.18 42.75 508.44 44.46 ;
   RECT 23.18 44.46 508.44 46.17 ;
   RECT 23.18 46.17 508.44 47.88 ;
   RECT 23.18 47.88 508.44 49.59 ;
   RECT 23.18 49.59 508.44 51.3 ;
   RECT 23.18 51.3 508.44 53.01 ;
   RECT 23.18 53.01 508.44 54.72 ;
   RECT 23.18 54.72 508.44 56.43 ;
   RECT 23.18 56.43 508.44 58.14 ;
   RECT 23.18 58.14 508.44 59.85 ;
   RECT 23.18 59.85 508.44 61.56 ;
   RECT 23.18 61.56 508.44 63.27 ;
   RECT 23.18 63.27 508.44 64.98 ;
   RECT 23.18 64.98 508.44 66.69 ;
   RECT 23.18 66.69 508.44 68.4 ;
   RECT 23.18 68.4 508.44 70.11 ;
   RECT 23.18 70.11 508.44 71.82 ;
   RECT 23.18 71.82 508.44 73.53 ;
   RECT 23.18 73.53 508.44 75.24 ;
   RECT 23.18 75.24 508.44 76.95 ;
   RECT 23.18 76.95 508.44 78.66 ;
   RECT 23.18 78.66 508.44 80.37 ;
   RECT 23.18 80.37 508.44 82.08 ;
   RECT 23.18 82.08 508.44 83.79 ;
   RECT 23.18 83.79 508.44 85.5 ;
   RECT 23.18 85.5 508.44 87.21 ;
   RECT 23.18 87.21 508.44 88.92 ;
   RECT 23.18 88.92 508.44 90.63 ;
   RECT 23.18 90.63 508.44 92.34 ;
   RECT 23.18 92.34 508.44 94.05 ;
   RECT 23.18 94.05 508.44 95.76 ;
   RECT 23.18 95.76 508.44 97.47 ;
   RECT 23.18 97.47 508.44 99.18 ;
   RECT 23.18 99.18 508.44 100.89 ;
   RECT 23.18 100.89 508.44 102.6 ;
   RECT 23.18 102.6 508.44 104.31 ;
   RECT 23.18 104.31 508.44 106.02 ;
   RECT 23.18 106.02 508.44 107.73 ;
   RECT 23.18 107.73 508.44 109.44 ;
   RECT 23.18 109.44 508.44 111.15 ;
   RECT 23.18 111.15 508.44 112.86 ;
   RECT 23.18 112.86 508.44 114.57 ;
   RECT 23.18 114.57 508.44 116.28 ;
   RECT 23.18 116.28 508.44 117.99 ;
   RECT 23.18 117.99 508.44 119.7 ;
   RECT 23.18 119.7 508.44 121.41 ;
   RECT 23.18 121.41 508.44 123.12 ;
   RECT 23.18 123.12 508.44 124.83 ;
   RECT 23.18 124.83 508.44 126.54 ;
   RECT 23.18 126.54 508.44 128.25 ;
   RECT 23.18 128.25 508.44 129.96 ;
   RECT 23.18 129.96 508.44 131.67 ;
   RECT 23.18 131.67 508.44 133.38 ;
   RECT 23.18 133.38 508.44 135.09 ;
   RECT 23.18 135.09 508.44 136.8 ;
   RECT 23.18 136.8 508.44 138.51 ;
   RECT 23.18 138.51 508.44 140.22 ;
   RECT 23.18 140.22 508.44 141.93 ;
   RECT 23.18 141.93 508.44 143.64 ;
   RECT 23.18 143.64 508.44 145.35 ;
   RECT 23.18 145.35 508.44 147.06 ;
   RECT 23.18 147.06 508.44 148.77 ;
   RECT 23.18 148.77 508.44 150.48 ;
   RECT 23.18 150.48 508.44 152.19 ;
   RECT 23.18 152.19 508.44 153.9 ;
   RECT 23.18 153.9 508.44 155.61 ;
   RECT 23.18 155.61 508.44 157.32 ;
   RECT 23.18 157.32 508.44 159.03 ;
   RECT 23.18 159.03 508.44 160.74 ;
   RECT 23.18 160.74 508.44 162.45 ;
   RECT 23.18 162.45 508.44 164.16 ;
   RECT 23.18 164.16 508.44 165.87 ;
   RECT 23.18 165.87 508.44 167.58 ;
   RECT 23.18 167.58 508.44 169.29 ;
   RECT 23.18 169.29 508.44 171.0 ;
   RECT 23.18 171.0 508.44 172.71 ;
   RECT 23.18 172.71 508.44 174.42 ;
   RECT 23.18 174.42 508.44 176.13 ;
   RECT 23.18 176.13 508.44 177.84 ;
   RECT 23.18 177.84 508.44 179.55 ;
   RECT 23.18 179.55 508.44 181.26 ;
   RECT 23.18 181.26 508.44 182.97 ;
   RECT 0.0 182.97 508.44 184.68 ;
   RECT 0.0 184.68 508.44 186.39 ;
   RECT 0.0 186.39 508.44 188.1 ;
   RECT 0.0 188.1 508.44 189.81 ;
   RECT 0.0 189.81 508.44 191.52 ;
   RECT 0.0 191.52 508.44 193.23 ;
   RECT 0.0 193.23 508.44 194.94 ;
   RECT 0.0 194.94 508.44 196.65 ;
   RECT 0.0 196.65 508.44 198.36 ;
   RECT 0.0 198.36 508.44 200.07 ;
   RECT 0.0 200.07 508.44 201.78 ;
   RECT 0.0 201.78 508.44 203.49 ;
   RECT 0.0 203.49 508.44 205.2 ;
   RECT 0.0 205.2 508.44 206.91 ;
   RECT 0.0 206.91 508.44 208.62 ;
   RECT 0.0 208.62 508.44 210.33 ;
   RECT 0.0 210.33 508.44 212.04 ;
   RECT 23.18 212.04 508.44 213.75 ;
   RECT 23.18 213.75 508.44 215.46 ;
   RECT 23.18 215.46 508.44 217.17 ;
   RECT 23.18 217.17 508.44 218.88 ;
   RECT 23.18 218.88 508.44 220.59 ;
   RECT 23.18 220.59 508.44 222.3 ;
   RECT 23.18 222.3 508.44 224.01 ;
   RECT 23.18 224.01 508.44 225.72 ;
   RECT 23.18 225.72 508.44 227.43 ;
   RECT 23.18 227.43 508.44 229.14 ;
   RECT 23.18 229.14 508.44 230.85 ;
   RECT 23.18 230.85 508.44 232.56 ;
   RECT 23.18 232.56 508.44 234.27 ;
   RECT 23.18 234.27 508.44 235.98 ;
   RECT 23.18 235.98 508.44 237.69 ;
   RECT 23.18 237.69 508.44 239.4 ;
   RECT 23.18 239.4 508.44 241.11 ;
   RECT 23.18 241.11 508.44 242.82 ;
   RECT 23.18 242.82 508.44 244.53 ;
   RECT 23.18 244.53 508.44 246.24 ;
   RECT 23.18 246.24 508.44 247.95 ;
   RECT 23.18 247.95 508.44 249.66 ;
   RECT 23.18 249.66 508.44 251.37 ;
   RECT 23.18 251.37 508.44 253.08 ;
   RECT 23.18 253.08 508.44 254.79 ;
   RECT 23.18 254.79 508.44 256.5 ;
   RECT 23.18 256.5 508.44 258.21 ;
   RECT 23.18 258.21 508.44 259.92 ;
   RECT 23.18 259.92 508.44 261.63 ;
   RECT 23.18 261.63 508.44 263.34 ;
   RECT 23.18 263.34 508.44 265.05 ;
   RECT 23.18 265.05 508.44 266.76 ;
   RECT 23.18 266.76 508.44 268.47 ;
   RECT 23.18 268.47 508.44 270.18 ;
   RECT 23.18 270.18 508.44 271.89 ;
   RECT 23.18 271.89 508.44 273.6 ;
   RECT 23.18 273.6 508.44 275.31 ;
   RECT 23.18 275.31 508.44 277.02 ;
   RECT 23.18 277.02 508.44 278.73 ;
   RECT 23.18 278.73 508.44 280.44 ;
   RECT 23.18 280.44 508.44 282.15 ;
   RECT 23.18 282.15 508.44 283.86 ;
   RECT 23.18 283.86 508.44 285.57 ;
   RECT 23.18 285.57 508.44 287.28 ;
   RECT 23.18 287.28 508.44 288.99 ;
   RECT 23.18 288.99 508.44 290.7 ;
   RECT 23.18 290.7 508.44 292.41 ;
   RECT 23.18 292.41 508.44 294.12 ;
   RECT 23.18 294.12 508.44 295.83 ;
   RECT 23.18 295.83 508.44 297.54 ;
   RECT 23.18 297.54 508.44 299.25 ;
   RECT 23.18 299.25 508.44 300.96 ;
   RECT 23.18 300.96 508.44 302.67 ;
   RECT 23.18 302.67 508.44 304.38 ;
   RECT 23.18 304.38 508.44 306.09 ;
   RECT 23.18 306.09 508.44 307.8 ;
   RECT 23.18 307.8 508.44 309.51 ;
   RECT 23.18 309.51 508.44 311.22 ;
   RECT 23.18 311.22 508.44 312.93 ;
   RECT 23.18 312.93 508.44 314.64 ;
   RECT 23.18 314.64 508.44 316.35 ;
   RECT 23.18 316.35 508.44 318.06 ;
   RECT 23.18 318.06 508.44 319.77 ;
   RECT 23.18 319.77 508.44 321.48 ;
   RECT 23.18 321.48 508.44 323.19 ;
   RECT 23.18 323.19 508.44 324.9 ;
   RECT 23.18 324.9 508.44 326.61 ;
   RECT 23.18 326.61 508.44 328.32 ;
   RECT 23.18 328.32 508.44 330.03 ;
   RECT 23.18 330.03 508.44 331.74 ;
   RECT 23.18 331.74 508.44 333.45 ;
   RECT 23.18 333.45 508.44 335.16 ;
   RECT 23.18 335.16 508.44 336.87 ;
   RECT 23.18 336.87 508.44 338.58 ;
   RECT 23.18 338.58 508.44 340.29 ;
   RECT 23.18 340.29 508.44 342.0 ;
   RECT 23.18 342.0 508.44 343.71 ;
   RECT 23.18 343.71 508.44 345.42 ;
   RECT 23.18 345.42 508.44 347.13 ;
   RECT 23.18 347.13 508.44 348.84 ;
   RECT 23.18 348.84 508.44 350.55 ;
   RECT 23.18 350.55 508.44 352.26 ;
   RECT 23.18 352.26 508.44 353.97 ;
   RECT 23.18 353.97 508.44 355.68 ;
   RECT 23.18 355.68 508.44 357.39 ;
   RECT 23.18 357.39 508.44 359.1 ;
   RECT 23.18 359.1 508.44 360.81 ;
   RECT 23.18 360.81 508.44 362.52 ;
   RECT 23.18 362.52 508.44 364.23 ;
   RECT 23.18 364.23 508.44 365.94 ;
   RECT 23.18 365.94 508.44 367.65 ;
   RECT 23.18 367.65 508.44 369.36 ;
   RECT 23.18 369.36 508.44 371.07 ;
   RECT 23.18 371.07 508.44 372.78 ;
   RECT 23.18 372.78 508.44 374.49 ;
   RECT 23.18 374.49 508.44 376.2 ;
   RECT 23.18 376.2 508.44 377.91 ;
   RECT 23.18 377.91 508.44 379.62 ;
   RECT 23.18 379.62 508.44 381.33 ;
   RECT 23.18 381.33 508.44 383.04 ;
   RECT 23.18 383.04 508.44 384.75 ;
   RECT 23.18 384.75 508.44 386.46 ;
   RECT 23.18 386.46 508.44 388.17 ;
   RECT 23.18 388.17 508.44 389.88 ;
   RECT 23.18 389.88 508.44 391.59 ;
   RECT 23.18 391.59 508.44 393.3 ;
   RECT 23.18 393.3 508.44 395.01 ;
   RECT 23.18 395.01 508.44 396.72 ;
   RECT 23.18 396.72 508.44 398.43 ;
   RECT 23.18 398.43 508.44 400.14 ;
   RECT 23.18 400.14 508.44 401.85 ;
   RECT 23.18 401.85 508.44 403.56 ;
   RECT 23.18 403.56 508.44 405.27 ;
   RECT 23.18 405.27 508.44 406.98 ;
   RECT 23.18 406.98 508.44 408.69 ;
   RECT 23.18 408.69 508.44 410.4 ;
 END
END block_1338x2160_145

MACRO block_533x1125_122
 CLASS BLOCK ;
 FOREIGN block_533x1125_122 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 202.54 BY 213.75 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 208.145 176.225 208.715 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 199.975 176.225 200.545 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 79.895 176.225 80.465 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 71.725 176.225 72.295 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 63.555 176.225 64.125 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 55.385 176.225 55.955 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 28.975 176.225 29.545 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 20.805 176.225 21.375 ;
  END
 END o7
 PIN o8
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 12.635 176.225 13.205 ;
  END
 END o8
 PIN o9
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 4.465 176.225 5.035 ;
  END
 END o9
 PIN o10
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 191.805 176.225 192.375 ;
  END
 END o10
 PIN o11
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 183.635 176.225 184.205 ;
  END
 END o11
 PIN o12
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 175.465 176.225 176.035 ;
  END
 END o12
 PIN o13
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 149.055 176.225 149.625 ;
  END
 END o13
 PIN o14
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 140.885 176.225 141.455 ;
  END
 END o14
 PIN o15
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 132.715 176.225 133.285 ;
  END
 END o15
 PIN o16
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 124.545 176.225 125.115 ;
  END
 END o16
 PIN o17
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 116.375 176.225 116.945 ;
  END
 END o17
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.835 109.345 199.405 109.915 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.835 92.245 199.405 92.815 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.835 104.025 199.405 104.595 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.835 99.655 199.405 100.225 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.075 108.965 198.645 109.535 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.075 109.725 198.645 110.295 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.835 110.105 199.405 110.675 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.835 100.415 199.405 100.985 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.835 87.305 199.405 87.875 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.075 92.625 198.645 93.195 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.835 93.005 199.405 93.575 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.835 90.915 199.405 91.485 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.835 88.445 199.405 89.015 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.075 86.925 198.645 87.495 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 188.955 110.485 189.525 111.055 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 188.955 97.185 189.525 97.755 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 209.855 176.225 210.425 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 201.685 176.225 202.255 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 78.185 176.225 78.755 ;
  END
 END i18
 PIN i19
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 70.015 176.225 70.585 ;
  END
 END i19
 PIN i20
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 61.845 176.225 62.415 ;
  END
 END i20
 PIN i21
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 53.675 176.225 54.245 ;
  END
 END i21
 PIN i22
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 27.265 176.225 27.835 ;
  END
 END i22
 PIN i23
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 19.095 176.225 19.665 ;
  END
 END i23
 PIN i24
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 10.925 176.225 11.495 ;
  END
 END i24
 PIN i25
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 2.755 176.225 3.325 ;
  END
 END i25
 PIN i26
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 193.515 176.225 194.085 ;
  END
 END i26
 PIN i27
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 185.345 176.225 185.915 ;
  END
 END i27
 PIN i28
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 177.175 176.225 177.745 ;
  END
 END i28
 PIN i29
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 150.765 176.225 151.335 ;
  END
 END i29
 PIN i30
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 142.595 176.225 143.165 ;
  END
 END i30
 PIN i31
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 134.425 176.225 134.995 ;
  END
 END i31
 PIN i32
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 126.255 176.225 126.825 ;
  END
 END i32
 PIN i33
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 118.085 176.225 118.655 ;
  END
 END i33
 PIN i34
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 195.225 176.225 195.795 ;
  END
 END i34
 PIN i35
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 191.235 175.465 191.805 ;
  END
 END i35
 PIN i36
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 187.055 176.225 187.625 ;
  END
 END i36
 PIN i37
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 203.395 176.225 203.965 ;
  END
 END i37
 PIN i38
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 127.965 176.225 128.535 ;
  END
 END i38
 PIN i39
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 123.975 175.465 124.545 ;
  END
 END i39
 PIN i40
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 119.795 176.225 120.365 ;
  END
 END i40
 PIN i41
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 115.805 175.465 116.375 ;
  END
 END i41
 PIN i42
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 76.475 176.225 77.045 ;
  END
 END i42
 PIN i43
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 80.465 175.465 81.035 ;
  END
 END i43
 PIN i44
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 84.645 176.225 85.215 ;
  END
 END i44
 PIN i45
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 68.305 176.225 68.875 ;
  END
 END i45
 PIN i46
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 9.215 176.225 9.785 ;
  END
 END i46
 PIN i47
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 13.205 175.465 13.775 ;
  END
 END i47
 PIN i48
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 17.385 176.225 17.955 ;
  END
 END i48
 PIN i49
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 21.375 175.465 21.945 ;
  END
 END i49
 PIN i50
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 199.405 175.465 199.975 ;
  END
 END i50
 PIN i51
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 132.145 175.465 132.715 ;
  END
 END i51
 PIN i52
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 72.295 175.465 72.865 ;
  END
 END i52
 PIN i53
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 5.035 175.465 5.605 ;
  END
 END i53
 PIN i54
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 184.015 110.485 184.585 111.055 ;
  END
 END i54
 PIN i55
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 184.015 97.185 184.585 97.755 ;
  END
 END i55
 PIN i56
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 209.285 175.465 209.855 ;
  END
 END i56
 PIN i57
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 201.115 175.465 201.685 ;
  END
 END i57
 PIN i58
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 78.755 175.465 79.325 ;
  END
 END i58
 PIN i59
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 70.585 175.465 71.155 ;
  END
 END i59
 PIN i60
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 62.415 175.465 62.985 ;
  END
 END i60
 PIN i61
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 54.245 175.465 54.815 ;
  END
 END i61
 PIN i62
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 27.835 175.465 28.405 ;
  END
 END i62
 PIN i63
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 19.665 175.465 20.235 ;
  END
 END i63
 PIN i64
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 11.495 175.465 12.065 ;
  END
 END i64
 PIN i65
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 3.325 175.465 3.895 ;
  END
 END i65
 PIN i66
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 192.945 175.465 193.515 ;
  END
 END i66
 PIN i67
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 184.775 175.465 185.345 ;
  END
 END i67
 PIN i68
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 176.605 175.465 177.175 ;
  END
 END i68
 PIN i69
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 150.195 175.465 150.765 ;
  END
 END i69
 PIN i70
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 142.025 175.465 142.595 ;
  END
 END i70
 PIN i71
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 133.855 175.465 134.425 ;
  END
 END i71
 PIN i72
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 125.685 175.465 126.255 ;
  END
 END i72
 PIN i73
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 117.515 175.465 118.085 ;
  END
 END i73
 PIN i74
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.835 102.885 199.405 103.455 ;
  END
 END i74
 PIN i75
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.075 102.505 198.645 103.075 ;
  END
 END i75
 PIN i76
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 208.715 174.705 209.285 ;
  END
 END i76
 PIN i77
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 200.545 174.705 201.115 ;
  END
 END i77
 PIN i78
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 79.325 174.705 79.895 ;
  END
 END i78
 PIN i79
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 71.155 174.705 71.725 ;
  END
 END i79
 PIN i80
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 62.985 174.705 63.555 ;
  END
 END i80
 PIN i81
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 54.815 174.705 55.385 ;
  END
 END i81
 PIN i82
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 28.405 174.705 28.975 ;
  END
 END i82
 PIN i83
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 20.235 174.705 20.805 ;
  END
 END i83
 PIN i84
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 12.065 174.705 12.635 ;
  END
 END i84
 PIN i85
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 3.895 174.705 4.465 ;
  END
 END i85
 PIN i86
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 192.375 174.705 192.945 ;
  END
 END i86
 PIN i87
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 184.205 174.705 184.775 ;
  END
 END i87
 PIN i88
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 176.035 174.705 176.605 ;
  END
 END i88
 PIN i89
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 149.625 174.705 150.195 ;
  END
 END i89
 PIN i90
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 141.455 174.705 142.025 ;
  END
 END i90
 PIN i91
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 133.285 174.705 133.855 ;
  END
 END i91
 PIN i92
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 125.115 174.705 125.685 ;
  END
 END i92
 PIN i93
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.135 116.945 174.705 117.515 ;
  END
 END i93
 PIN i94
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 197.695 110.485 198.265 111.055 ;
  END
 END i94
 PIN i95
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 196.555 110.485 197.125 111.055 ;
  END
 END i95
 PIN i96
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 195.035 110.485 195.605 111.055 ;
  END
 END i96
 PIN i97
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 193.135 110.485 193.705 111.055 ;
  END
 END i97
 PIN i98
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 191.995 110.485 192.565 111.055 ;
  END
 END i98
 PIN i99
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 197.695 97.185 198.265 97.755 ;
  END
 END i99
 PIN i100
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 196.555 97.185 197.125 97.755 ;
  END
 END i100
 PIN i101
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 195.035 97.185 195.605 97.755 ;
  END
 END i101
 PIN i102
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 193.135 97.185 193.705 97.755 ;
  END
 END i102
 PIN i103
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 191.995 97.185 192.565 97.755 ;
  END
 END i103
 OBS
  LAYER metal1 ;
   RECT 0.0 0.0 179.36 1.71 ;
   RECT 0.0 1.71 179.36 3.42 ;
   RECT 0.0 3.42 179.36 5.13 ;
   RECT 0.0 5.13 179.36 6.84 ;
   RECT 0.0 6.84 179.36 8.55 ;
   RECT 0.0 8.55 179.36 10.26 ;
   RECT 0.0 10.26 179.36 11.97 ;
   RECT 0.0 11.97 179.36 13.68 ;
   RECT 0.0 13.68 179.36 15.39 ;
   RECT 0.0 15.39 179.36 17.1 ;
   RECT 0.0 17.1 179.36 18.81 ;
   RECT 0.0 18.81 179.36 20.52 ;
   RECT 0.0 20.52 179.36 22.23 ;
   RECT 0.0 22.23 179.36 23.94 ;
   RECT 0.0 23.94 179.36 25.65 ;
   RECT 0.0 25.65 179.36 27.36 ;
   RECT 0.0 27.36 179.36 29.07 ;
   RECT 0.0 29.07 179.36 30.78 ;
   RECT 0.0 30.78 179.36 32.49 ;
   RECT 0.0 32.49 179.36 34.2 ;
   RECT 0.0 34.2 179.36 35.91 ;
   RECT 0.0 35.91 179.36 37.62 ;
   RECT 0.0 37.62 179.36 39.33 ;
   RECT 0.0 39.33 179.36 41.04 ;
   RECT 0.0 41.04 179.36 42.75 ;
   RECT 0.0 42.75 179.36 44.46 ;
   RECT 0.0 44.46 179.36 46.17 ;
   RECT 0.0 46.17 179.36 47.88 ;
   RECT 0.0 47.88 179.36 49.59 ;
   RECT 0.0 49.59 179.36 51.3 ;
   RECT 0.0 51.3 179.36 53.01 ;
   RECT 0.0 53.01 179.36 54.72 ;
   RECT 0.0 54.72 179.36 56.43 ;
   RECT 0.0 56.43 179.36 58.14 ;
   RECT 0.0 58.14 179.36 59.85 ;
   RECT 0.0 59.85 179.36 61.56 ;
   RECT 0.0 61.56 179.36 63.27 ;
   RECT 0.0 63.27 179.36 64.98 ;
   RECT 0.0 64.98 179.36 66.69 ;
   RECT 0.0 66.69 179.36 68.4 ;
   RECT 0.0 68.4 179.36 70.11 ;
   RECT 0.0 70.11 179.36 71.82 ;
   RECT 0.0 71.82 179.36 73.53 ;
   RECT 0.0 73.53 179.36 75.24 ;
   RECT 0.0 75.24 179.36 76.95 ;
   RECT 0.0 76.95 179.36 78.66 ;
   RECT 0.0 78.66 179.36 80.37 ;
   RECT 0.0 80.37 179.36 82.08 ;
   RECT 0.0 82.08 179.36 83.79 ;
   RECT 0.0 83.79 202.54 85.5 ;
   RECT 0.0 85.5 202.54 87.21 ;
   RECT 0.0 87.21 202.54 88.92 ;
   RECT 0.0 88.92 202.54 90.63 ;
   RECT 0.0 90.63 202.54 92.34 ;
   RECT 0.0 92.34 202.54 94.05 ;
   RECT 0.0 94.05 202.54 95.76 ;
   RECT 0.0 95.76 202.54 97.47 ;
   RECT 0.0 97.47 202.54 99.18 ;
   RECT 0.0 99.18 202.54 100.89 ;
   RECT 0.0 100.89 202.54 102.6 ;
   RECT 0.0 102.6 202.54 104.31 ;
   RECT 0.0 104.31 202.54 106.02 ;
   RECT 0.0 106.02 202.54 107.73 ;
   RECT 0.0 107.73 202.54 109.44 ;
   RECT 0.0 109.44 202.54 111.15 ;
   RECT 0.0 111.15 202.54 112.86 ;
   RECT 0.0 112.86 179.36 114.57 ;
   RECT 0.0 114.57 179.36 116.28 ;
   RECT 0.0 116.28 179.36 117.99 ;
   RECT 0.0 117.99 179.36 119.7 ;
   RECT 0.0 119.7 179.36 121.41 ;
   RECT 0.0 121.41 179.36 123.12 ;
   RECT 0.0 123.12 179.36 124.83 ;
   RECT 0.0 124.83 179.36 126.54 ;
   RECT 0.0 126.54 179.36 128.25 ;
   RECT 0.0 128.25 179.36 129.96 ;
   RECT 0.0 129.96 179.36 131.67 ;
   RECT 0.0 131.67 179.36 133.38 ;
   RECT 0.0 133.38 179.36 135.09 ;
   RECT 0.0 135.09 179.36 136.8 ;
   RECT 0.0 136.8 179.36 138.51 ;
   RECT 0.0 138.51 179.36 140.22 ;
   RECT 0.0 140.22 179.36 141.93 ;
   RECT 0.0 141.93 179.36 143.64 ;
   RECT 0.0 143.64 179.36 145.35 ;
   RECT 0.0 145.35 179.36 147.06 ;
   RECT 0.0 147.06 179.36 148.77 ;
   RECT 0.0 148.77 179.36 150.48 ;
   RECT 0.0 150.48 179.36 152.19 ;
   RECT 0.0 152.19 179.36 153.9 ;
   RECT 0.0 153.9 179.36 155.61 ;
   RECT 0.0 155.61 179.36 157.32 ;
   RECT 0.0 157.32 179.36 159.03 ;
   RECT 0.0 159.03 179.36 160.74 ;
   RECT 0.0 160.74 179.36 162.45 ;
   RECT 0.0 162.45 179.36 164.16 ;
   RECT 0.0 164.16 179.36 165.87 ;
   RECT 0.0 165.87 179.36 167.58 ;
   RECT 0.0 167.58 179.36 169.29 ;
   RECT 0.0 169.29 179.36 171.0 ;
   RECT 0.0 171.0 179.36 172.71 ;
   RECT 0.0 172.71 179.36 174.42 ;
   RECT 0.0 174.42 179.36 176.13 ;
   RECT 0.0 176.13 179.36 177.84 ;
   RECT 0.0 177.84 179.36 179.55 ;
   RECT 0.0 179.55 179.36 181.26 ;
   RECT 0.0 181.26 179.36 182.97 ;
   RECT 0.0 182.97 179.36 184.68 ;
   RECT 0.0 184.68 179.36 186.39 ;
   RECT 0.0 186.39 179.36 188.1 ;
   RECT 0.0 188.1 179.36 189.81 ;
   RECT 0.0 189.81 179.36 191.52 ;
   RECT 0.0 191.52 179.36 193.23 ;
   RECT 0.0 193.23 179.36 194.94 ;
   RECT 0.0 194.94 179.36 196.65 ;
   RECT 0.0 196.65 179.36 198.36 ;
   RECT 0.0 198.36 179.36 200.07 ;
   RECT 0.0 200.07 179.36 201.78 ;
   RECT 0.0 201.78 179.36 203.49 ;
   RECT 0.0 203.49 179.36 205.2 ;
   RECT 0.0 205.2 179.36 206.91 ;
   RECT 0.0 206.91 179.36 208.62 ;
   RECT 0.0 208.62 179.36 210.33 ;
   RECT 0.0 210.33 179.36 212.04 ;
   RECT 0.0 212.04 179.36 213.75 ;
  LAYER via1 ;
   RECT 0.0 0.0 179.36 1.71 ;
   RECT 0.0 1.71 179.36 3.42 ;
   RECT 0.0 3.42 179.36 5.13 ;
   RECT 0.0 5.13 179.36 6.84 ;
   RECT 0.0 6.84 179.36 8.55 ;
   RECT 0.0 8.55 179.36 10.26 ;
   RECT 0.0 10.26 179.36 11.97 ;
   RECT 0.0 11.97 179.36 13.68 ;
   RECT 0.0 13.68 179.36 15.39 ;
   RECT 0.0 15.39 179.36 17.1 ;
   RECT 0.0 17.1 179.36 18.81 ;
   RECT 0.0 18.81 179.36 20.52 ;
   RECT 0.0 20.52 179.36 22.23 ;
   RECT 0.0 22.23 179.36 23.94 ;
   RECT 0.0 23.94 179.36 25.65 ;
   RECT 0.0 25.65 179.36 27.36 ;
   RECT 0.0 27.36 179.36 29.07 ;
   RECT 0.0 29.07 179.36 30.78 ;
   RECT 0.0 30.78 179.36 32.49 ;
   RECT 0.0 32.49 179.36 34.2 ;
   RECT 0.0 34.2 179.36 35.91 ;
   RECT 0.0 35.91 179.36 37.62 ;
   RECT 0.0 37.62 179.36 39.33 ;
   RECT 0.0 39.33 179.36 41.04 ;
   RECT 0.0 41.04 179.36 42.75 ;
   RECT 0.0 42.75 179.36 44.46 ;
   RECT 0.0 44.46 179.36 46.17 ;
   RECT 0.0 46.17 179.36 47.88 ;
   RECT 0.0 47.88 179.36 49.59 ;
   RECT 0.0 49.59 179.36 51.3 ;
   RECT 0.0 51.3 179.36 53.01 ;
   RECT 0.0 53.01 179.36 54.72 ;
   RECT 0.0 54.72 179.36 56.43 ;
   RECT 0.0 56.43 179.36 58.14 ;
   RECT 0.0 58.14 179.36 59.85 ;
   RECT 0.0 59.85 179.36 61.56 ;
   RECT 0.0 61.56 179.36 63.27 ;
   RECT 0.0 63.27 179.36 64.98 ;
   RECT 0.0 64.98 179.36 66.69 ;
   RECT 0.0 66.69 179.36 68.4 ;
   RECT 0.0 68.4 179.36 70.11 ;
   RECT 0.0 70.11 179.36 71.82 ;
   RECT 0.0 71.82 179.36 73.53 ;
   RECT 0.0 73.53 179.36 75.24 ;
   RECT 0.0 75.24 179.36 76.95 ;
   RECT 0.0 76.95 179.36 78.66 ;
   RECT 0.0 78.66 179.36 80.37 ;
   RECT 0.0 80.37 179.36 82.08 ;
   RECT 0.0 82.08 179.36 83.79 ;
   RECT 0.0 83.79 202.54 85.5 ;
   RECT 0.0 85.5 202.54 87.21 ;
   RECT 0.0 87.21 202.54 88.92 ;
   RECT 0.0 88.92 202.54 90.63 ;
   RECT 0.0 90.63 202.54 92.34 ;
   RECT 0.0 92.34 202.54 94.05 ;
   RECT 0.0 94.05 202.54 95.76 ;
   RECT 0.0 95.76 202.54 97.47 ;
   RECT 0.0 97.47 202.54 99.18 ;
   RECT 0.0 99.18 202.54 100.89 ;
   RECT 0.0 100.89 202.54 102.6 ;
   RECT 0.0 102.6 202.54 104.31 ;
   RECT 0.0 104.31 202.54 106.02 ;
   RECT 0.0 106.02 202.54 107.73 ;
   RECT 0.0 107.73 202.54 109.44 ;
   RECT 0.0 109.44 202.54 111.15 ;
   RECT 0.0 111.15 202.54 112.86 ;
   RECT 0.0 112.86 179.36 114.57 ;
   RECT 0.0 114.57 179.36 116.28 ;
   RECT 0.0 116.28 179.36 117.99 ;
   RECT 0.0 117.99 179.36 119.7 ;
   RECT 0.0 119.7 179.36 121.41 ;
   RECT 0.0 121.41 179.36 123.12 ;
   RECT 0.0 123.12 179.36 124.83 ;
   RECT 0.0 124.83 179.36 126.54 ;
   RECT 0.0 126.54 179.36 128.25 ;
   RECT 0.0 128.25 179.36 129.96 ;
   RECT 0.0 129.96 179.36 131.67 ;
   RECT 0.0 131.67 179.36 133.38 ;
   RECT 0.0 133.38 179.36 135.09 ;
   RECT 0.0 135.09 179.36 136.8 ;
   RECT 0.0 136.8 179.36 138.51 ;
   RECT 0.0 138.51 179.36 140.22 ;
   RECT 0.0 140.22 179.36 141.93 ;
   RECT 0.0 141.93 179.36 143.64 ;
   RECT 0.0 143.64 179.36 145.35 ;
   RECT 0.0 145.35 179.36 147.06 ;
   RECT 0.0 147.06 179.36 148.77 ;
   RECT 0.0 148.77 179.36 150.48 ;
   RECT 0.0 150.48 179.36 152.19 ;
   RECT 0.0 152.19 179.36 153.9 ;
   RECT 0.0 153.9 179.36 155.61 ;
   RECT 0.0 155.61 179.36 157.32 ;
   RECT 0.0 157.32 179.36 159.03 ;
   RECT 0.0 159.03 179.36 160.74 ;
   RECT 0.0 160.74 179.36 162.45 ;
   RECT 0.0 162.45 179.36 164.16 ;
   RECT 0.0 164.16 179.36 165.87 ;
   RECT 0.0 165.87 179.36 167.58 ;
   RECT 0.0 167.58 179.36 169.29 ;
   RECT 0.0 169.29 179.36 171.0 ;
   RECT 0.0 171.0 179.36 172.71 ;
   RECT 0.0 172.71 179.36 174.42 ;
   RECT 0.0 174.42 179.36 176.13 ;
   RECT 0.0 176.13 179.36 177.84 ;
   RECT 0.0 177.84 179.36 179.55 ;
   RECT 0.0 179.55 179.36 181.26 ;
   RECT 0.0 181.26 179.36 182.97 ;
   RECT 0.0 182.97 179.36 184.68 ;
   RECT 0.0 184.68 179.36 186.39 ;
   RECT 0.0 186.39 179.36 188.1 ;
   RECT 0.0 188.1 179.36 189.81 ;
   RECT 0.0 189.81 179.36 191.52 ;
   RECT 0.0 191.52 179.36 193.23 ;
   RECT 0.0 193.23 179.36 194.94 ;
   RECT 0.0 194.94 179.36 196.65 ;
   RECT 0.0 196.65 179.36 198.36 ;
   RECT 0.0 198.36 179.36 200.07 ;
   RECT 0.0 200.07 179.36 201.78 ;
   RECT 0.0 201.78 179.36 203.49 ;
   RECT 0.0 203.49 179.36 205.2 ;
   RECT 0.0 205.2 179.36 206.91 ;
   RECT 0.0 206.91 179.36 208.62 ;
   RECT 0.0 208.62 179.36 210.33 ;
   RECT 0.0 210.33 179.36 212.04 ;
   RECT 0.0 212.04 179.36 213.75 ;
  LAYER metal2 ;
   RECT 0.0 0.0 179.36 1.71 ;
   RECT 0.0 1.71 179.36 3.42 ;
   RECT 0.0 3.42 179.36 5.13 ;
   RECT 0.0 5.13 179.36 6.84 ;
   RECT 0.0 6.84 179.36 8.55 ;
   RECT 0.0 8.55 179.36 10.26 ;
   RECT 0.0 10.26 179.36 11.97 ;
   RECT 0.0 11.97 179.36 13.68 ;
   RECT 0.0 13.68 179.36 15.39 ;
   RECT 0.0 15.39 179.36 17.1 ;
   RECT 0.0 17.1 179.36 18.81 ;
   RECT 0.0 18.81 179.36 20.52 ;
   RECT 0.0 20.52 179.36 22.23 ;
   RECT 0.0 22.23 179.36 23.94 ;
   RECT 0.0 23.94 179.36 25.65 ;
   RECT 0.0 25.65 179.36 27.36 ;
   RECT 0.0 27.36 179.36 29.07 ;
   RECT 0.0 29.07 179.36 30.78 ;
   RECT 0.0 30.78 179.36 32.49 ;
   RECT 0.0 32.49 179.36 34.2 ;
   RECT 0.0 34.2 179.36 35.91 ;
   RECT 0.0 35.91 179.36 37.62 ;
   RECT 0.0 37.62 179.36 39.33 ;
   RECT 0.0 39.33 179.36 41.04 ;
   RECT 0.0 41.04 179.36 42.75 ;
   RECT 0.0 42.75 179.36 44.46 ;
   RECT 0.0 44.46 179.36 46.17 ;
   RECT 0.0 46.17 179.36 47.88 ;
   RECT 0.0 47.88 179.36 49.59 ;
   RECT 0.0 49.59 179.36 51.3 ;
   RECT 0.0 51.3 179.36 53.01 ;
   RECT 0.0 53.01 179.36 54.72 ;
   RECT 0.0 54.72 179.36 56.43 ;
   RECT 0.0 56.43 179.36 58.14 ;
   RECT 0.0 58.14 179.36 59.85 ;
   RECT 0.0 59.85 179.36 61.56 ;
   RECT 0.0 61.56 179.36 63.27 ;
   RECT 0.0 63.27 179.36 64.98 ;
   RECT 0.0 64.98 179.36 66.69 ;
   RECT 0.0 66.69 179.36 68.4 ;
   RECT 0.0 68.4 179.36 70.11 ;
   RECT 0.0 70.11 179.36 71.82 ;
   RECT 0.0 71.82 179.36 73.53 ;
   RECT 0.0 73.53 179.36 75.24 ;
   RECT 0.0 75.24 179.36 76.95 ;
   RECT 0.0 76.95 179.36 78.66 ;
   RECT 0.0 78.66 179.36 80.37 ;
   RECT 0.0 80.37 179.36 82.08 ;
   RECT 0.0 82.08 179.36 83.79 ;
   RECT 0.0 83.79 202.54 85.5 ;
   RECT 0.0 85.5 202.54 87.21 ;
   RECT 0.0 87.21 202.54 88.92 ;
   RECT 0.0 88.92 202.54 90.63 ;
   RECT 0.0 90.63 202.54 92.34 ;
   RECT 0.0 92.34 202.54 94.05 ;
   RECT 0.0 94.05 202.54 95.76 ;
   RECT 0.0 95.76 202.54 97.47 ;
   RECT 0.0 97.47 202.54 99.18 ;
   RECT 0.0 99.18 202.54 100.89 ;
   RECT 0.0 100.89 202.54 102.6 ;
   RECT 0.0 102.6 202.54 104.31 ;
   RECT 0.0 104.31 202.54 106.02 ;
   RECT 0.0 106.02 202.54 107.73 ;
   RECT 0.0 107.73 202.54 109.44 ;
   RECT 0.0 109.44 202.54 111.15 ;
   RECT 0.0 111.15 202.54 112.86 ;
   RECT 0.0 112.86 179.36 114.57 ;
   RECT 0.0 114.57 179.36 116.28 ;
   RECT 0.0 116.28 179.36 117.99 ;
   RECT 0.0 117.99 179.36 119.7 ;
   RECT 0.0 119.7 179.36 121.41 ;
   RECT 0.0 121.41 179.36 123.12 ;
   RECT 0.0 123.12 179.36 124.83 ;
   RECT 0.0 124.83 179.36 126.54 ;
   RECT 0.0 126.54 179.36 128.25 ;
   RECT 0.0 128.25 179.36 129.96 ;
   RECT 0.0 129.96 179.36 131.67 ;
   RECT 0.0 131.67 179.36 133.38 ;
   RECT 0.0 133.38 179.36 135.09 ;
   RECT 0.0 135.09 179.36 136.8 ;
   RECT 0.0 136.8 179.36 138.51 ;
   RECT 0.0 138.51 179.36 140.22 ;
   RECT 0.0 140.22 179.36 141.93 ;
   RECT 0.0 141.93 179.36 143.64 ;
   RECT 0.0 143.64 179.36 145.35 ;
   RECT 0.0 145.35 179.36 147.06 ;
   RECT 0.0 147.06 179.36 148.77 ;
   RECT 0.0 148.77 179.36 150.48 ;
   RECT 0.0 150.48 179.36 152.19 ;
   RECT 0.0 152.19 179.36 153.9 ;
   RECT 0.0 153.9 179.36 155.61 ;
   RECT 0.0 155.61 179.36 157.32 ;
   RECT 0.0 157.32 179.36 159.03 ;
   RECT 0.0 159.03 179.36 160.74 ;
   RECT 0.0 160.74 179.36 162.45 ;
   RECT 0.0 162.45 179.36 164.16 ;
   RECT 0.0 164.16 179.36 165.87 ;
   RECT 0.0 165.87 179.36 167.58 ;
   RECT 0.0 167.58 179.36 169.29 ;
   RECT 0.0 169.29 179.36 171.0 ;
   RECT 0.0 171.0 179.36 172.71 ;
   RECT 0.0 172.71 179.36 174.42 ;
   RECT 0.0 174.42 179.36 176.13 ;
   RECT 0.0 176.13 179.36 177.84 ;
   RECT 0.0 177.84 179.36 179.55 ;
   RECT 0.0 179.55 179.36 181.26 ;
   RECT 0.0 181.26 179.36 182.97 ;
   RECT 0.0 182.97 179.36 184.68 ;
   RECT 0.0 184.68 179.36 186.39 ;
   RECT 0.0 186.39 179.36 188.1 ;
   RECT 0.0 188.1 179.36 189.81 ;
   RECT 0.0 189.81 179.36 191.52 ;
   RECT 0.0 191.52 179.36 193.23 ;
   RECT 0.0 193.23 179.36 194.94 ;
   RECT 0.0 194.94 179.36 196.65 ;
   RECT 0.0 196.65 179.36 198.36 ;
   RECT 0.0 198.36 179.36 200.07 ;
   RECT 0.0 200.07 179.36 201.78 ;
   RECT 0.0 201.78 179.36 203.49 ;
   RECT 0.0 203.49 179.36 205.2 ;
   RECT 0.0 205.2 179.36 206.91 ;
   RECT 0.0 206.91 179.36 208.62 ;
   RECT 0.0 208.62 179.36 210.33 ;
   RECT 0.0 210.33 179.36 212.04 ;
   RECT 0.0 212.04 179.36 213.75 ;
  LAYER via2 ;
   RECT 0.0 0.0 179.36 1.71 ;
   RECT 0.0 1.71 179.36 3.42 ;
   RECT 0.0 3.42 179.36 5.13 ;
   RECT 0.0 5.13 179.36 6.84 ;
   RECT 0.0 6.84 179.36 8.55 ;
   RECT 0.0 8.55 179.36 10.26 ;
   RECT 0.0 10.26 179.36 11.97 ;
   RECT 0.0 11.97 179.36 13.68 ;
   RECT 0.0 13.68 179.36 15.39 ;
   RECT 0.0 15.39 179.36 17.1 ;
   RECT 0.0 17.1 179.36 18.81 ;
   RECT 0.0 18.81 179.36 20.52 ;
   RECT 0.0 20.52 179.36 22.23 ;
   RECT 0.0 22.23 179.36 23.94 ;
   RECT 0.0 23.94 179.36 25.65 ;
   RECT 0.0 25.65 179.36 27.36 ;
   RECT 0.0 27.36 179.36 29.07 ;
   RECT 0.0 29.07 179.36 30.78 ;
   RECT 0.0 30.78 179.36 32.49 ;
   RECT 0.0 32.49 179.36 34.2 ;
   RECT 0.0 34.2 179.36 35.91 ;
   RECT 0.0 35.91 179.36 37.62 ;
   RECT 0.0 37.62 179.36 39.33 ;
   RECT 0.0 39.33 179.36 41.04 ;
   RECT 0.0 41.04 179.36 42.75 ;
   RECT 0.0 42.75 179.36 44.46 ;
   RECT 0.0 44.46 179.36 46.17 ;
   RECT 0.0 46.17 179.36 47.88 ;
   RECT 0.0 47.88 179.36 49.59 ;
   RECT 0.0 49.59 179.36 51.3 ;
   RECT 0.0 51.3 179.36 53.01 ;
   RECT 0.0 53.01 179.36 54.72 ;
   RECT 0.0 54.72 179.36 56.43 ;
   RECT 0.0 56.43 179.36 58.14 ;
   RECT 0.0 58.14 179.36 59.85 ;
   RECT 0.0 59.85 179.36 61.56 ;
   RECT 0.0 61.56 179.36 63.27 ;
   RECT 0.0 63.27 179.36 64.98 ;
   RECT 0.0 64.98 179.36 66.69 ;
   RECT 0.0 66.69 179.36 68.4 ;
   RECT 0.0 68.4 179.36 70.11 ;
   RECT 0.0 70.11 179.36 71.82 ;
   RECT 0.0 71.82 179.36 73.53 ;
   RECT 0.0 73.53 179.36 75.24 ;
   RECT 0.0 75.24 179.36 76.95 ;
   RECT 0.0 76.95 179.36 78.66 ;
   RECT 0.0 78.66 179.36 80.37 ;
   RECT 0.0 80.37 179.36 82.08 ;
   RECT 0.0 82.08 179.36 83.79 ;
   RECT 0.0 83.79 202.54 85.5 ;
   RECT 0.0 85.5 202.54 87.21 ;
   RECT 0.0 87.21 202.54 88.92 ;
   RECT 0.0 88.92 202.54 90.63 ;
   RECT 0.0 90.63 202.54 92.34 ;
   RECT 0.0 92.34 202.54 94.05 ;
   RECT 0.0 94.05 202.54 95.76 ;
   RECT 0.0 95.76 202.54 97.47 ;
   RECT 0.0 97.47 202.54 99.18 ;
   RECT 0.0 99.18 202.54 100.89 ;
   RECT 0.0 100.89 202.54 102.6 ;
   RECT 0.0 102.6 202.54 104.31 ;
   RECT 0.0 104.31 202.54 106.02 ;
   RECT 0.0 106.02 202.54 107.73 ;
   RECT 0.0 107.73 202.54 109.44 ;
   RECT 0.0 109.44 202.54 111.15 ;
   RECT 0.0 111.15 202.54 112.86 ;
   RECT 0.0 112.86 179.36 114.57 ;
   RECT 0.0 114.57 179.36 116.28 ;
   RECT 0.0 116.28 179.36 117.99 ;
   RECT 0.0 117.99 179.36 119.7 ;
   RECT 0.0 119.7 179.36 121.41 ;
   RECT 0.0 121.41 179.36 123.12 ;
   RECT 0.0 123.12 179.36 124.83 ;
   RECT 0.0 124.83 179.36 126.54 ;
   RECT 0.0 126.54 179.36 128.25 ;
   RECT 0.0 128.25 179.36 129.96 ;
   RECT 0.0 129.96 179.36 131.67 ;
   RECT 0.0 131.67 179.36 133.38 ;
   RECT 0.0 133.38 179.36 135.09 ;
   RECT 0.0 135.09 179.36 136.8 ;
   RECT 0.0 136.8 179.36 138.51 ;
   RECT 0.0 138.51 179.36 140.22 ;
   RECT 0.0 140.22 179.36 141.93 ;
   RECT 0.0 141.93 179.36 143.64 ;
   RECT 0.0 143.64 179.36 145.35 ;
   RECT 0.0 145.35 179.36 147.06 ;
   RECT 0.0 147.06 179.36 148.77 ;
   RECT 0.0 148.77 179.36 150.48 ;
   RECT 0.0 150.48 179.36 152.19 ;
   RECT 0.0 152.19 179.36 153.9 ;
   RECT 0.0 153.9 179.36 155.61 ;
   RECT 0.0 155.61 179.36 157.32 ;
   RECT 0.0 157.32 179.36 159.03 ;
   RECT 0.0 159.03 179.36 160.74 ;
   RECT 0.0 160.74 179.36 162.45 ;
   RECT 0.0 162.45 179.36 164.16 ;
   RECT 0.0 164.16 179.36 165.87 ;
   RECT 0.0 165.87 179.36 167.58 ;
   RECT 0.0 167.58 179.36 169.29 ;
   RECT 0.0 169.29 179.36 171.0 ;
   RECT 0.0 171.0 179.36 172.71 ;
   RECT 0.0 172.71 179.36 174.42 ;
   RECT 0.0 174.42 179.36 176.13 ;
   RECT 0.0 176.13 179.36 177.84 ;
   RECT 0.0 177.84 179.36 179.55 ;
   RECT 0.0 179.55 179.36 181.26 ;
   RECT 0.0 181.26 179.36 182.97 ;
   RECT 0.0 182.97 179.36 184.68 ;
   RECT 0.0 184.68 179.36 186.39 ;
   RECT 0.0 186.39 179.36 188.1 ;
   RECT 0.0 188.1 179.36 189.81 ;
   RECT 0.0 189.81 179.36 191.52 ;
   RECT 0.0 191.52 179.36 193.23 ;
   RECT 0.0 193.23 179.36 194.94 ;
   RECT 0.0 194.94 179.36 196.65 ;
   RECT 0.0 196.65 179.36 198.36 ;
   RECT 0.0 198.36 179.36 200.07 ;
   RECT 0.0 200.07 179.36 201.78 ;
   RECT 0.0 201.78 179.36 203.49 ;
   RECT 0.0 203.49 179.36 205.2 ;
   RECT 0.0 205.2 179.36 206.91 ;
   RECT 0.0 206.91 179.36 208.62 ;
   RECT 0.0 208.62 179.36 210.33 ;
   RECT 0.0 210.33 179.36 212.04 ;
   RECT 0.0 212.04 179.36 213.75 ;
  LAYER metal3 ;
   RECT 0.0 0.0 179.36 1.71 ;
   RECT 0.0 1.71 179.36 3.42 ;
   RECT 0.0 3.42 179.36 5.13 ;
   RECT 0.0 5.13 179.36 6.84 ;
   RECT 0.0 6.84 179.36 8.55 ;
   RECT 0.0 8.55 179.36 10.26 ;
   RECT 0.0 10.26 179.36 11.97 ;
   RECT 0.0 11.97 179.36 13.68 ;
   RECT 0.0 13.68 179.36 15.39 ;
   RECT 0.0 15.39 179.36 17.1 ;
   RECT 0.0 17.1 179.36 18.81 ;
   RECT 0.0 18.81 179.36 20.52 ;
   RECT 0.0 20.52 179.36 22.23 ;
   RECT 0.0 22.23 179.36 23.94 ;
   RECT 0.0 23.94 179.36 25.65 ;
   RECT 0.0 25.65 179.36 27.36 ;
   RECT 0.0 27.36 179.36 29.07 ;
   RECT 0.0 29.07 179.36 30.78 ;
   RECT 0.0 30.78 179.36 32.49 ;
   RECT 0.0 32.49 179.36 34.2 ;
   RECT 0.0 34.2 179.36 35.91 ;
   RECT 0.0 35.91 179.36 37.62 ;
   RECT 0.0 37.62 179.36 39.33 ;
   RECT 0.0 39.33 179.36 41.04 ;
   RECT 0.0 41.04 179.36 42.75 ;
   RECT 0.0 42.75 179.36 44.46 ;
   RECT 0.0 44.46 179.36 46.17 ;
   RECT 0.0 46.17 179.36 47.88 ;
   RECT 0.0 47.88 179.36 49.59 ;
   RECT 0.0 49.59 179.36 51.3 ;
   RECT 0.0 51.3 179.36 53.01 ;
   RECT 0.0 53.01 179.36 54.72 ;
   RECT 0.0 54.72 179.36 56.43 ;
   RECT 0.0 56.43 179.36 58.14 ;
   RECT 0.0 58.14 179.36 59.85 ;
   RECT 0.0 59.85 179.36 61.56 ;
   RECT 0.0 61.56 179.36 63.27 ;
   RECT 0.0 63.27 179.36 64.98 ;
   RECT 0.0 64.98 179.36 66.69 ;
   RECT 0.0 66.69 179.36 68.4 ;
   RECT 0.0 68.4 179.36 70.11 ;
   RECT 0.0 70.11 179.36 71.82 ;
   RECT 0.0 71.82 179.36 73.53 ;
   RECT 0.0 73.53 179.36 75.24 ;
   RECT 0.0 75.24 179.36 76.95 ;
   RECT 0.0 76.95 179.36 78.66 ;
   RECT 0.0 78.66 179.36 80.37 ;
   RECT 0.0 80.37 179.36 82.08 ;
   RECT 0.0 82.08 179.36 83.79 ;
   RECT 0.0 83.79 202.54 85.5 ;
   RECT 0.0 85.5 202.54 87.21 ;
   RECT 0.0 87.21 202.54 88.92 ;
   RECT 0.0 88.92 202.54 90.63 ;
   RECT 0.0 90.63 202.54 92.34 ;
   RECT 0.0 92.34 202.54 94.05 ;
   RECT 0.0 94.05 202.54 95.76 ;
   RECT 0.0 95.76 202.54 97.47 ;
   RECT 0.0 97.47 202.54 99.18 ;
   RECT 0.0 99.18 202.54 100.89 ;
   RECT 0.0 100.89 202.54 102.6 ;
   RECT 0.0 102.6 202.54 104.31 ;
   RECT 0.0 104.31 202.54 106.02 ;
   RECT 0.0 106.02 202.54 107.73 ;
   RECT 0.0 107.73 202.54 109.44 ;
   RECT 0.0 109.44 202.54 111.15 ;
   RECT 0.0 111.15 202.54 112.86 ;
   RECT 0.0 112.86 179.36 114.57 ;
   RECT 0.0 114.57 179.36 116.28 ;
   RECT 0.0 116.28 179.36 117.99 ;
   RECT 0.0 117.99 179.36 119.7 ;
   RECT 0.0 119.7 179.36 121.41 ;
   RECT 0.0 121.41 179.36 123.12 ;
   RECT 0.0 123.12 179.36 124.83 ;
   RECT 0.0 124.83 179.36 126.54 ;
   RECT 0.0 126.54 179.36 128.25 ;
   RECT 0.0 128.25 179.36 129.96 ;
   RECT 0.0 129.96 179.36 131.67 ;
   RECT 0.0 131.67 179.36 133.38 ;
   RECT 0.0 133.38 179.36 135.09 ;
   RECT 0.0 135.09 179.36 136.8 ;
   RECT 0.0 136.8 179.36 138.51 ;
   RECT 0.0 138.51 179.36 140.22 ;
   RECT 0.0 140.22 179.36 141.93 ;
   RECT 0.0 141.93 179.36 143.64 ;
   RECT 0.0 143.64 179.36 145.35 ;
   RECT 0.0 145.35 179.36 147.06 ;
   RECT 0.0 147.06 179.36 148.77 ;
   RECT 0.0 148.77 179.36 150.48 ;
   RECT 0.0 150.48 179.36 152.19 ;
   RECT 0.0 152.19 179.36 153.9 ;
   RECT 0.0 153.9 179.36 155.61 ;
   RECT 0.0 155.61 179.36 157.32 ;
   RECT 0.0 157.32 179.36 159.03 ;
   RECT 0.0 159.03 179.36 160.74 ;
   RECT 0.0 160.74 179.36 162.45 ;
   RECT 0.0 162.45 179.36 164.16 ;
   RECT 0.0 164.16 179.36 165.87 ;
   RECT 0.0 165.87 179.36 167.58 ;
   RECT 0.0 167.58 179.36 169.29 ;
   RECT 0.0 169.29 179.36 171.0 ;
   RECT 0.0 171.0 179.36 172.71 ;
   RECT 0.0 172.71 179.36 174.42 ;
   RECT 0.0 174.42 179.36 176.13 ;
   RECT 0.0 176.13 179.36 177.84 ;
   RECT 0.0 177.84 179.36 179.55 ;
   RECT 0.0 179.55 179.36 181.26 ;
   RECT 0.0 181.26 179.36 182.97 ;
   RECT 0.0 182.97 179.36 184.68 ;
   RECT 0.0 184.68 179.36 186.39 ;
   RECT 0.0 186.39 179.36 188.1 ;
   RECT 0.0 188.1 179.36 189.81 ;
   RECT 0.0 189.81 179.36 191.52 ;
   RECT 0.0 191.52 179.36 193.23 ;
   RECT 0.0 193.23 179.36 194.94 ;
   RECT 0.0 194.94 179.36 196.65 ;
   RECT 0.0 196.65 179.36 198.36 ;
   RECT 0.0 198.36 179.36 200.07 ;
   RECT 0.0 200.07 179.36 201.78 ;
   RECT 0.0 201.78 179.36 203.49 ;
   RECT 0.0 203.49 179.36 205.2 ;
   RECT 0.0 205.2 179.36 206.91 ;
   RECT 0.0 206.91 179.36 208.62 ;
   RECT 0.0 208.62 179.36 210.33 ;
   RECT 0.0 210.33 179.36 212.04 ;
   RECT 0.0 212.04 179.36 213.75 ;
  LAYER via3 ;
   RECT 0.0 0.0 179.36 1.71 ;
   RECT 0.0 1.71 179.36 3.42 ;
   RECT 0.0 3.42 179.36 5.13 ;
   RECT 0.0 5.13 179.36 6.84 ;
   RECT 0.0 6.84 179.36 8.55 ;
   RECT 0.0 8.55 179.36 10.26 ;
   RECT 0.0 10.26 179.36 11.97 ;
   RECT 0.0 11.97 179.36 13.68 ;
   RECT 0.0 13.68 179.36 15.39 ;
   RECT 0.0 15.39 179.36 17.1 ;
   RECT 0.0 17.1 179.36 18.81 ;
   RECT 0.0 18.81 179.36 20.52 ;
   RECT 0.0 20.52 179.36 22.23 ;
   RECT 0.0 22.23 179.36 23.94 ;
   RECT 0.0 23.94 179.36 25.65 ;
   RECT 0.0 25.65 179.36 27.36 ;
   RECT 0.0 27.36 179.36 29.07 ;
   RECT 0.0 29.07 179.36 30.78 ;
   RECT 0.0 30.78 179.36 32.49 ;
   RECT 0.0 32.49 179.36 34.2 ;
   RECT 0.0 34.2 179.36 35.91 ;
   RECT 0.0 35.91 179.36 37.62 ;
   RECT 0.0 37.62 179.36 39.33 ;
   RECT 0.0 39.33 179.36 41.04 ;
   RECT 0.0 41.04 179.36 42.75 ;
   RECT 0.0 42.75 179.36 44.46 ;
   RECT 0.0 44.46 179.36 46.17 ;
   RECT 0.0 46.17 179.36 47.88 ;
   RECT 0.0 47.88 179.36 49.59 ;
   RECT 0.0 49.59 179.36 51.3 ;
   RECT 0.0 51.3 179.36 53.01 ;
   RECT 0.0 53.01 179.36 54.72 ;
   RECT 0.0 54.72 179.36 56.43 ;
   RECT 0.0 56.43 179.36 58.14 ;
   RECT 0.0 58.14 179.36 59.85 ;
   RECT 0.0 59.85 179.36 61.56 ;
   RECT 0.0 61.56 179.36 63.27 ;
   RECT 0.0 63.27 179.36 64.98 ;
   RECT 0.0 64.98 179.36 66.69 ;
   RECT 0.0 66.69 179.36 68.4 ;
   RECT 0.0 68.4 179.36 70.11 ;
   RECT 0.0 70.11 179.36 71.82 ;
   RECT 0.0 71.82 179.36 73.53 ;
   RECT 0.0 73.53 179.36 75.24 ;
   RECT 0.0 75.24 179.36 76.95 ;
   RECT 0.0 76.95 179.36 78.66 ;
   RECT 0.0 78.66 179.36 80.37 ;
   RECT 0.0 80.37 179.36 82.08 ;
   RECT 0.0 82.08 179.36 83.79 ;
   RECT 0.0 83.79 202.54 85.5 ;
   RECT 0.0 85.5 202.54 87.21 ;
   RECT 0.0 87.21 202.54 88.92 ;
   RECT 0.0 88.92 202.54 90.63 ;
   RECT 0.0 90.63 202.54 92.34 ;
   RECT 0.0 92.34 202.54 94.05 ;
   RECT 0.0 94.05 202.54 95.76 ;
   RECT 0.0 95.76 202.54 97.47 ;
   RECT 0.0 97.47 202.54 99.18 ;
   RECT 0.0 99.18 202.54 100.89 ;
   RECT 0.0 100.89 202.54 102.6 ;
   RECT 0.0 102.6 202.54 104.31 ;
   RECT 0.0 104.31 202.54 106.02 ;
   RECT 0.0 106.02 202.54 107.73 ;
   RECT 0.0 107.73 202.54 109.44 ;
   RECT 0.0 109.44 202.54 111.15 ;
   RECT 0.0 111.15 202.54 112.86 ;
   RECT 0.0 112.86 179.36 114.57 ;
   RECT 0.0 114.57 179.36 116.28 ;
   RECT 0.0 116.28 179.36 117.99 ;
   RECT 0.0 117.99 179.36 119.7 ;
   RECT 0.0 119.7 179.36 121.41 ;
   RECT 0.0 121.41 179.36 123.12 ;
   RECT 0.0 123.12 179.36 124.83 ;
   RECT 0.0 124.83 179.36 126.54 ;
   RECT 0.0 126.54 179.36 128.25 ;
   RECT 0.0 128.25 179.36 129.96 ;
   RECT 0.0 129.96 179.36 131.67 ;
   RECT 0.0 131.67 179.36 133.38 ;
   RECT 0.0 133.38 179.36 135.09 ;
   RECT 0.0 135.09 179.36 136.8 ;
   RECT 0.0 136.8 179.36 138.51 ;
   RECT 0.0 138.51 179.36 140.22 ;
   RECT 0.0 140.22 179.36 141.93 ;
   RECT 0.0 141.93 179.36 143.64 ;
   RECT 0.0 143.64 179.36 145.35 ;
   RECT 0.0 145.35 179.36 147.06 ;
   RECT 0.0 147.06 179.36 148.77 ;
   RECT 0.0 148.77 179.36 150.48 ;
   RECT 0.0 150.48 179.36 152.19 ;
   RECT 0.0 152.19 179.36 153.9 ;
   RECT 0.0 153.9 179.36 155.61 ;
   RECT 0.0 155.61 179.36 157.32 ;
   RECT 0.0 157.32 179.36 159.03 ;
   RECT 0.0 159.03 179.36 160.74 ;
   RECT 0.0 160.74 179.36 162.45 ;
   RECT 0.0 162.45 179.36 164.16 ;
   RECT 0.0 164.16 179.36 165.87 ;
   RECT 0.0 165.87 179.36 167.58 ;
   RECT 0.0 167.58 179.36 169.29 ;
   RECT 0.0 169.29 179.36 171.0 ;
   RECT 0.0 171.0 179.36 172.71 ;
   RECT 0.0 172.71 179.36 174.42 ;
   RECT 0.0 174.42 179.36 176.13 ;
   RECT 0.0 176.13 179.36 177.84 ;
   RECT 0.0 177.84 179.36 179.55 ;
   RECT 0.0 179.55 179.36 181.26 ;
   RECT 0.0 181.26 179.36 182.97 ;
   RECT 0.0 182.97 179.36 184.68 ;
   RECT 0.0 184.68 179.36 186.39 ;
   RECT 0.0 186.39 179.36 188.1 ;
   RECT 0.0 188.1 179.36 189.81 ;
   RECT 0.0 189.81 179.36 191.52 ;
   RECT 0.0 191.52 179.36 193.23 ;
   RECT 0.0 193.23 179.36 194.94 ;
   RECT 0.0 194.94 179.36 196.65 ;
   RECT 0.0 196.65 179.36 198.36 ;
   RECT 0.0 198.36 179.36 200.07 ;
   RECT 0.0 200.07 179.36 201.78 ;
   RECT 0.0 201.78 179.36 203.49 ;
   RECT 0.0 203.49 179.36 205.2 ;
   RECT 0.0 205.2 179.36 206.91 ;
   RECT 0.0 206.91 179.36 208.62 ;
   RECT 0.0 208.62 179.36 210.33 ;
   RECT 0.0 210.33 179.36 212.04 ;
   RECT 0.0 212.04 179.36 213.75 ;
  LAYER metal4 ;
   RECT 0.0 0.0 179.36 1.71 ;
   RECT 0.0 1.71 179.36 3.42 ;
   RECT 0.0 3.42 179.36 5.13 ;
   RECT 0.0 5.13 179.36 6.84 ;
   RECT 0.0 6.84 179.36 8.55 ;
   RECT 0.0 8.55 179.36 10.26 ;
   RECT 0.0 10.26 179.36 11.97 ;
   RECT 0.0 11.97 179.36 13.68 ;
   RECT 0.0 13.68 179.36 15.39 ;
   RECT 0.0 15.39 179.36 17.1 ;
   RECT 0.0 17.1 179.36 18.81 ;
   RECT 0.0 18.81 179.36 20.52 ;
   RECT 0.0 20.52 179.36 22.23 ;
   RECT 0.0 22.23 179.36 23.94 ;
   RECT 0.0 23.94 179.36 25.65 ;
   RECT 0.0 25.65 179.36 27.36 ;
   RECT 0.0 27.36 179.36 29.07 ;
   RECT 0.0 29.07 179.36 30.78 ;
   RECT 0.0 30.78 179.36 32.49 ;
   RECT 0.0 32.49 179.36 34.2 ;
   RECT 0.0 34.2 179.36 35.91 ;
   RECT 0.0 35.91 179.36 37.62 ;
   RECT 0.0 37.62 179.36 39.33 ;
   RECT 0.0 39.33 179.36 41.04 ;
   RECT 0.0 41.04 179.36 42.75 ;
   RECT 0.0 42.75 179.36 44.46 ;
   RECT 0.0 44.46 179.36 46.17 ;
   RECT 0.0 46.17 179.36 47.88 ;
   RECT 0.0 47.88 179.36 49.59 ;
   RECT 0.0 49.59 179.36 51.3 ;
   RECT 0.0 51.3 179.36 53.01 ;
   RECT 0.0 53.01 179.36 54.72 ;
   RECT 0.0 54.72 179.36 56.43 ;
   RECT 0.0 56.43 179.36 58.14 ;
   RECT 0.0 58.14 179.36 59.85 ;
   RECT 0.0 59.85 179.36 61.56 ;
   RECT 0.0 61.56 179.36 63.27 ;
   RECT 0.0 63.27 179.36 64.98 ;
   RECT 0.0 64.98 179.36 66.69 ;
   RECT 0.0 66.69 179.36 68.4 ;
   RECT 0.0 68.4 179.36 70.11 ;
   RECT 0.0 70.11 179.36 71.82 ;
   RECT 0.0 71.82 179.36 73.53 ;
   RECT 0.0 73.53 179.36 75.24 ;
   RECT 0.0 75.24 179.36 76.95 ;
   RECT 0.0 76.95 179.36 78.66 ;
   RECT 0.0 78.66 179.36 80.37 ;
   RECT 0.0 80.37 179.36 82.08 ;
   RECT 0.0 82.08 179.36 83.79 ;
   RECT 0.0 83.79 202.54 85.5 ;
   RECT 0.0 85.5 202.54 87.21 ;
   RECT 0.0 87.21 202.54 88.92 ;
   RECT 0.0 88.92 202.54 90.63 ;
   RECT 0.0 90.63 202.54 92.34 ;
   RECT 0.0 92.34 202.54 94.05 ;
   RECT 0.0 94.05 202.54 95.76 ;
   RECT 0.0 95.76 202.54 97.47 ;
   RECT 0.0 97.47 202.54 99.18 ;
   RECT 0.0 99.18 202.54 100.89 ;
   RECT 0.0 100.89 202.54 102.6 ;
   RECT 0.0 102.6 202.54 104.31 ;
   RECT 0.0 104.31 202.54 106.02 ;
   RECT 0.0 106.02 202.54 107.73 ;
   RECT 0.0 107.73 202.54 109.44 ;
   RECT 0.0 109.44 202.54 111.15 ;
   RECT 0.0 111.15 202.54 112.86 ;
   RECT 0.0 112.86 179.36 114.57 ;
   RECT 0.0 114.57 179.36 116.28 ;
   RECT 0.0 116.28 179.36 117.99 ;
   RECT 0.0 117.99 179.36 119.7 ;
   RECT 0.0 119.7 179.36 121.41 ;
   RECT 0.0 121.41 179.36 123.12 ;
   RECT 0.0 123.12 179.36 124.83 ;
   RECT 0.0 124.83 179.36 126.54 ;
   RECT 0.0 126.54 179.36 128.25 ;
   RECT 0.0 128.25 179.36 129.96 ;
   RECT 0.0 129.96 179.36 131.67 ;
   RECT 0.0 131.67 179.36 133.38 ;
   RECT 0.0 133.38 179.36 135.09 ;
   RECT 0.0 135.09 179.36 136.8 ;
   RECT 0.0 136.8 179.36 138.51 ;
   RECT 0.0 138.51 179.36 140.22 ;
   RECT 0.0 140.22 179.36 141.93 ;
   RECT 0.0 141.93 179.36 143.64 ;
   RECT 0.0 143.64 179.36 145.35 ;
   RECT 0.0 145.35 179.36 147.06 ;
   RECT 0.0 147.06 179.36 148.77 ;
   RECT 0.0 148.77 179.36 150.48 ;
   RECT 0.0 150.48 179.36 152.19 ;
   RECT 0.0 152.19 179.36 153.9 ;
   RECT 0.0 153.9 179.36 155.61 ;
   RECT 0.0 155.61 179.36 157.32 ;
   RECT 0.0 157.32 179.36 159.03 ;
   RECT 0.0 159.03 179.36 160.74 ;
   RECT 0.0 160.74 179.36 162.45 ;
   RECT 0.0 162.45 179.36 164.16 ;
   RECT 0.0 164.16 179.36 165.87 ;
   RECT 0.0 165.87 179.36 167.58 ;
   RECT 0.0 167.58 179.36 169.29 ;
   RECT 0.0 169.29 179.36 171.0 ;
   RECT 0.0 171.0 179.36 172.71 ;
   RECT 0.0 172.71 179.36 174.42 ;
   RECT 0.0 174.42 179.36 176.13 ;
   RECT 0.0 176.13 179.36 177.84 ;
   RECT 0.0 177.84 179.36 179.55 ;
   RECT 0.0 179.55 179.36 181.26 ;
   RECT 0.0 181.26 179.36 182.97 ;
   RECT 0.0 182.97 179.36 184.68 ;
   RECT 0.0 184.68 179.36 186.39 ;
   RECT 0.0 186.39 179.36 188.1 ;
   RECT 0.0 188.1 179.36 189.81 ;
   RECT 0.0 189.81 179.36 191.52 ;
   RECT 0.0 191.52 179.36 193.23 ;
   RECT 0.0 193.23 179.36 194.94 ;
   RECT 0.0 194.94 179.36 196.65 ;
   RECT 0.0 196.65 179.36 198.36 ;
   RECT 0.0 198.36 179.36 200.07 ;
   RECT 0.0 200.07 179.36 201.78 ;
   RECT 0.0 201.78 179.36 203.49 ;
   RECT 0.0 203.49 179.36 205.2 ;
   RECT 0.0 205.2 179.36 206.91 ;
   RECT 0.0 206.91 179.36 208.62 ;
   RECT 0.0 208.62 179.36 210.33 ;
   RECT 0.0 210.33 179.36 212.04 ;
   RECT 0.0 212.04 179.36 213.75 ;
 END
END block_533x1125_122

MACRO block_1829x2160_148
 CLASS BLOCK ;
 FOREIGN block_1829x2160_148 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 695.02 BY 410.4 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 400.045 668.705 400.615 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 383.705 668.705 384.275 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 218.405 668.705 218.975 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 173.945 668.705 174.515 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 157.605 668.705 158.175 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 141.265 668.705 141.835 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 124.925 668.705 125.495 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 108.585 668.705 109.155 ;
  END
 END o7
 PIN o8
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 74.005 668.705 74.575 ;
  END
 END o8
 PIN o9
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 57.665 668.705 58.235 ;
  END
 END o9
 PIN o10
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 41.325 668.705 41.895 ;
  END
 END o10
 PIN o11
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 24.985 668.705 25.555 ;
  END
 END o11
 PIN o12
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 367.365 668.705 367.935 ;
  END
 END o12
 PIN o13
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 8.645 668.705 9.215 ;
  END
 END o13
 PIN o14
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 351.025 668.705 351.595 ;
  END
 END o14
 PIN o15
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 334.685 668.705 335.255 ;
  END
 END o15
 PIN o16
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 318.345 668.705 318.915 ;
  END
 END o16
 PIN o17
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 283.765 668.705 284.335 ;
  END
 END o17
 PIN o18
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 267.425 668.705 267.995 ;
  END
 END o18
 PIN o19
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 251.085 668.705 251.655 ;
  END
 END o19
 PIN o20
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 234.745 668.705 235.315 ;
  END
 END o20
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 691.315 207.385 691.885 207.955 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 691.315 185.725 691.885 186.295 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 691.315 190.285 691.885 190.855 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 691.315 202.065 691.885 202.635 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 691.315 197.695 691.885 198.265 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 691.315 194.845 691.885 195.415 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 690.555 207.005 691.125 207.575 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 690.555 207.765 691.125 208.335 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 691.315 208.145 691.885 208.715 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 691.315 198.455 691.885 199.025 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 690.555 185.345 691.125 185.915 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 690.555 190.665 691.125 191.235 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 691.315 193.895 691.885 194.465 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 691.315 186.485 691.885 187.055 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 691.315 191.045 691.885 191.615 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 691.315 188.955 691.885 189.525 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 690.555 186.105 691.125 186.675 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 691.315 184.965 691.885 185.535 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 680.295 208.525 680.865 209.095 ;
  END
 END i18
 PIN i19
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 678.395 208.525 678.965 209.095 ;
  END
 END i19
 PIN i20
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 680.295 195.225 680.865 195.795 ;
  END
 END i20
 PIN i21
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 678.395 195.225 678.965 195.795 ;
  END
 END i21
 PIN i22
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 401.755 668.705 402.325 ;
  END
 END i22
 PIN i23
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 385.415 668.705 385.985 ;
  END
 END i23
 PIN i24
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 220.115 668.705 220.685 ;
  END
 END i24
 PIN i25
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 172.235 668.705 172.805 ;
  END
 END i25
 PIN i26
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 155.895 668.705 156.465 ;
  END
 END i26
 PIN i27
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 139.555 668.705 140.125 ;
  END
 END i27
 PIN i28
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 123.215 668.705 123.785 ;
  END
 END i28
 PIN i29
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 106.875 668.705 107.445 ;
  END
 END i29
 PIN i30
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 72.295 668.705 72.865 ;
  END
 END i30
 PIN i31
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 55.955 668.705 56.525 ;
  END
 END i31
 PIN i32
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 39.615 668.705 40.185 ;
  END
 END i32
 PIN i33
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 23.275 668.705 23.845 ;
  END
 END i33
 PIN i34
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 369.075 668.705 369.645 ;
  END
 END i34
 PIN i35
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 6.935 668.705 7.505 ;
  END
 END i35
 PIN i36
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 352.735 668.705 353.305 ;
  END
 END i36
 PIN i37
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 336.395 668.705 336.965 ;
  END
 END i37
 PIN i38
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 320.055 668.705 320.625 ;
  END
 END i38
 PIN i39
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 285.475 668.705 286.045 ;
  END
 END i39
 PIN i40
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 269.135 668.705 269.705 ;
  END
 END i40
 PIN i41
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 252.795 668.705 253.365 ;
  END
 END i41
 PIN i42
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 236.455 668.705 237.025 ;
  END
 END i42
 PIN i43
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 667.375 334.115 667.945 334.685 ;
  END
 END i43
 PIN i44
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 330.125 668.705 330.695 ;
  END
 END i44
 PIN i45
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 325.945 668.705 326.515 ;
  END
 END i45
 PIN i46
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 346.465 668.705 347.035 ;
  END
 END i46
 PIN i47
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 342.285 668.705 342.855 ;
  END
 END i47
 PIN i48
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 667.375 266.855 667.945 267.425 ;
  END
 END i48
 PIN i49
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 262.865 668.705 263.435 ;
  END
 END i49
 PIN i50
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 258.685 668.705 259.255 ;
  END
 END i50
 PIN i51
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 254.695 668.705 255.265 ;
  END
 END i51
 PIN i52
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 667.375 250.515 667.945 251.085 ;
  END
 END i52
 PIN i53
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 667.375 125.495 667.945 126.065 ;
  END
 END i53
 PIN i54
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 129.485 668.705 130.055 ;
  END
 END i54
 PIN i55
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 133.665 668.705 134.235 ;
  END
 END i55
 PIN i56
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 137.655 668.705 138.225 ;
  END
 END i56
 PIN i57
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 667.375 141.835 667.945 142.405 ;
  END
 END i57
 PIN i58
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 667.375 58.235 667.945 58.805 ;
  END
 END i58
 PIN i59
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 62.225 668.705 62.795 ;
  END
 END i59
 PIN i60
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 66.405 668.705 66.975 ;
  END
 END i60
 PIN i61
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 45.885 668.705 46.455 ;
  END
 END i61
 PIN i62
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 50.065 668.705 50.635 ;
  END
 END i62
 PIN i63
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 338.295 668.705 338.865 ;
  END
 END i63
 PIN i64
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 271.035 668.705 271.605 ;
  END
 END i64
 PIN i65
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 121.315 668.705 121.885 ;
  END
 END i65
 PIN i66
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 668.135 54.055 668.705 54.625 ;
  END
 END i66
 PIN i67
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 676.495 208.525 677.065 209.095 ;
  END
 END i67
 PIN i68
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 676.495 195.225 677.065 195.795 ;
  END
 END i68
 PIN i69
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 667.375 401.185 667.945 401.755 ;
  END
 END i69
 PIN i70
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 667.375 384.845 667.945 385.415 ;
  END
 END i70
 PIN i71
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 667.375 219.545 667.945 220.115 ;
  END
 END i71
 PIN i72
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 667.375 172.805 667.945 173.375 ;
  END
 END i72
 PIN i73
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 667.375 156.465 667.945 157.035 ;
  END
 END i73
 PIN i74
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 667.375 140.125 667.945 140.695 ;
  END
 END i74
 PIN i75
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 667.375 123.785 667.945 124.355 ;
  END
 END i75
 PIN i76
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 667.375 107.445 667.945 108.015 ;
  END
 END i76
 PIN i77
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 667.375 72.865 667.945 73.435 ;
  END
 END i77
 PIN i78
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 667.375 56.525 667.945 57.095 ;
  END
 END i78
 PIN i79
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 667.375 40.185 667.945 40.755 ;
  END
 END i79
 PIN i80
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 667.375 23.845 667.945 24.415 ;
  END
 END i80
 PIN i81
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 667.375 368.505 667.945 369.075 ;
  END
 END i81
 PIN i82
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 667.375 7.505 667.945 8.075 ;
  END
 END i82
 PIN i83
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 667.375 352.165 667.945 352.735 ;
  END
 END i83
 PIN i84
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 667.375 335.825 667.945 336.395 ;
  END
 END i84
 PIN i85
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 667.375 319.485 667.945 320.055 ;
  END
 END i85
 PIN i86
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 667.375 284.905 667.945 285.475 ;
  END
 END i86
 PIN i87
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 667.375 268.565 667.945 269.135 ;
  END
 END i87
 PIN i88
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 667.375 252.225 667.945 252.795 ;
  END
 END i88
 PIN i89
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 667.375 235.885 667.945 236.455 ;
  END
 END i89
 PIN i90
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 691.315 200.925 691.885 201.495 ;
  END
 END i90
 PIN i91
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 690.555 200.545 691.125 201.115 ;
  END
 END i91
 PIN i92
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 666.615 400.615 667.185 401.185 ;
  END
 END i92
 PIN i93
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 666.615 384.275 667.185 384.845 ;
  END
 END i93
 PIN i94
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 666.615 218.975 667.185 219.545 ;
  END
 END i94
 PIN i95
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 666.615 173.375 667.185 173.945 ;
  END
 END i95
 PIN i96
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 666.615 157.035 667.185 157.605 ;
  END
 END i96
 PIN i97
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 666.615 140.695 667.185 141.265 ;
  END
 END i97
 PIN i98
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 666.615 124.355 667.185 124.925 ;
  END
 END i98
 PIN i99
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 666.615 108.015 667.185 108.585 ;
  END
 END i99
 PIN i100
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 666.615 73.435 667.185 74.005 ;
  END
 END i100
 PIN i101
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 666.615 57.095 667.185 57.665 ;
  END
 END i101
 PIN i102
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 666.615 40.755 667.185 41.325 ;
  END
 END i102
 PIN i103
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 666.615 24.415 667.185 24.985 ;
  END
 END i103
 PIN i104
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 666.615 367.935 667.185 368.505 ;
  END
 END i104
 PIN i105
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 666.615 8.075 667.185 8.645 ;
  END
 END i105
 PIN i106
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 666.615 351.595 667.185 352.165 ;
  END
 END i106
 PIN i107
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 666.615 335.255 667.185 335.825 ;
  END
 END i107
 PIN i108
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 666.615 318.915 667.185 319.485 ;
  END
 END i108
 PIN i109
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 666.615 284.335 667.185 284.905 ;
  END
 END i109
 PIN i110
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 666.615 267.995 667.185 268.565 ;
  END
 END i110
 PIN i111
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 666.615 251.655 667.185 252.225 ;
  END
 END i111
 PIN i112
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 666.615 235.315 667.185 235.885 ;
  END
 END i112
 PIN i113
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 690.175 208.525 690.745 209.095 ;
  END
 END i113
 PIN i114
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 689.035 208.525 689.605 209.095 ;
  END
 END i114
 PIN i115
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 687.515 208.525 688.085 209.095 ;
  END
 END i115
 PIN i116
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 685.615 208.525 686.185 209.095 ;
  END
 END i116
 PIN i117
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 684.095 208.525 684.665 209.095 ;
  END
 END i117
 PIN i118
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 682.575 208.525 683.145 209.095 ;
  END
 END i118
 PIN i119
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 681.435 208.525 682.005 209.095 ;
  END
 END i119
 PIN i120
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 690.175 195.225 690.745 195.795 ;
  END
 END i120
 PIN i121
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 689.035 195.225 689.605 195.795 ;
  END
 END i121
 PIN i122
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 687.515 195.225 688.085 195.795 ;
  END
 END i122
 PIN i123
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 685.615 195.225 686.185 195.795 ;
  END
 END i123
 PIN i124
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 684.095 195.225 684.665 195.795 ;
  END
 END i124
 PIN i125
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 682.575 195.225 683.145 195.795 ;
  END
 END i125
 PIN i126
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 681.435 195.225 682.005 195.795 ;
  END
 END i126
 OBS
  LAYER metal1 ;
   RECT 0.0 0.0 671.84 1.71 ;
   RECT 0.0 1.71 671.84 3.42 ;
   RECT 0.0 3.42 671.84 5.13 ;
   RECT 0.0 5.13 671.84 6.84 ;
   RECT 0.0 6.84 671.84 8.55 ;
   RECT 0.0 8.55 671.84 10.26 ;
   RECT 0.0 10.26 671.84 11.97 ;
   RECT 0.0 11.97 671.84 13.68 ;
   RECT 0.0 13.68 671.84 15.39 ;
   RECT 0.0 15.39 671.84 17.1 ;
   RECT 0.0 17.1 671.84 18.81 ;
   RECT 0.0 18.81 671.84 20.52 ;
   RECT 0.0 20.52 671.84 22.23 ;
   RECT 0.0 22.23 671.84 23.94 ;
   RECT 0.0 23.94 671.84 25.65 ;
   RECT 0.0 25.65 671.84 27.36 ;
   RECT 0.0 27.36 671.84 29.07 ;
   RECT 0.0 29.07 671.84 30.78 ;
   RECT 0.0 30.78 671.84 32.49 ;
   RECT 0.0 32.49 671.84 34.2 ;
   RECT 0.0 34.2 671.84 35.91 ;
   RECT 0.0 35.91 671.84 37.62 ;
   RECT 0.0 37.62 671.84 39.33 ;
   RECT 0.0 39.33 671.84 41.04 ;
   RECT 0.0 41.04 671.84 42.75 ;
   RECT 0.0 42.75 671.84 44.46 ;
   RECT 0.0 44.46 671.84 46.17 ;
   RECT 0.0 46.17 671.84 47.88 ;
   RECT 0.0 47.88 671.84 49.59 ;
   RECT 0.0 49.59 671.84 51.3 ;
   RECT 0.0 51.3 671.84 53.01 ;
   RECT 0.0 53.01 671.84 54.72 ;
   RECT 0.0 54.72 671.84 56.43 ;
   RECT 0.0 56.43 671.84 58.14 ;
   RECT 0.0 58.14 671.84 59.85 ;
   RECT 0.0 59.85 671.84 61.56 ;
   RECT 0.0 61.56 671.84 63.27 ;
   RECT 0.0 63.27 671.84 64.98 ;
   RECT 0.0 64.98 671.84 66.69 ;
   RECT 0.0 66.69 671.84 68.4 ;
   RECT 0.0 68.4 671.84 70.11 ;
   RECT 0.0 70.11 671.84 71.82 ;
   RECT 0.0 71.82 671.84 73.53 ;
   RECT 0.0 73.53 671.84 75.24 ;
   RECT 0.0 75.24 671.84 76.95 ;
   RECT 0.0 76.95 671.84 78.66 ;
   RECT 0.0 78.66 671.84 80.37 ;
   RECT 0.0 80.37 671.84 82.08 ;
   RECT 0.0 82.08 671.84 83.79 ;
   RECT 0.0 83.79 671.84 85.5 ;
   RECT 0.0 85.5 671.84 87.21 ;
   RECT 0.0 87.21 671.84 88.92 ;
   RECT 0.0 88.92 671.84 90.63 ;
   RECT 0.0 90.63 671.84 92.34 ;
   RECT 0.0 92.34 671.84 94.05 ;
   RECT 0.0 94.05 671.84 95.76 ;
   RECT 0.0 95.76 671.84 97.47 ;
   RECT 0.0 97.47 671.84 99.18 ;
   RECT 0.0 99.18 671.84 100.89 ;
   RECT 0.0 100.89 671.84 102.6 ;
   RECT 0.0 102.6 671.84 104.31 ;
   RECT 0.0 104.31 671.84 106.02 ;
   RECT 0.0 106.02 671.84 107.73 ;
   RECT 0.0 107.73 671.84 109.44 ;
   RECT 0.0 109.44 671.84 111.15 ;
   RECT 0.0 111.15 671.84 112.86 ;
   RECT 0.0 112.86 671.84 114.57 ;
   RECT 0.0 114.57 671.84 116.28 ;
   RECT 0.0 116.28 671.84 117.99 ;
   RECT 0.0 117.99 671.84 119.7 ;
   RECT 0.0 119.7 671.84 121.41 ;
   RECT 0.0 121.41 671.84 123.12 ;
   RECT 0.0 123.12 671.84 124.83 ;
   RECT 0.0 124.83 671.84 126.54 ;
   RECT 0.0 126.54 671.84 128.25 ;
   RECT 0.0 128.25 671.84 129.96 ;
   RECT 0.0 129.96 671.84 131.67 ;
   RECT 0.0 131.67 671.84 133.38 ;
   RECT 0.0 133.38 671.84 135.09 ;
   RECT 0.0 135.09 671.84 136.8 ;
   RECT 0.0 136.8 671.84 138.51 ;
   RECT 0.0 138.51 671.84 140.22 ;
   RECT 0.0 140.22 671.84 141.93 ;
   RECT 0.0 141.93 671.84 143.64 ;
   RECT 0.0 143.64 671.84 145.35 ;
   RECT 0.0 145.35 671.84 147.06 ;
   RECT 0.0 147.06 671.84 148.77 ;
   RECT 0.0 148.77 671.84 150.48 ;
   RECT 0.0 150.48 671.84 152.19 ;
   RECT 0.0 152.19 671.84 153.9 ;
   RECT 0.0 153.9 671.84 155.61 ;
   RECT 0.0 155.61 671.84 157.32 ;
   RECT 0.0 157.32 671.84 159.03 ;
   RECT 0.0 159.03 671.84 160.74 ;
   RECT 0.0 160.74 671.84 162.45 ;
   RECT 0.0 162.45 671.84 164.16 ;
   RECT 0.0 164.16 671.84 165.87 ;
   RECT 0.0 165.87 671.84 167.58 ;
   RECT 0.0 167.58 671.84 169.29 ;
   RECT 0.0 169.29 671.84 171.0 ;
   RECT 0.0 171.0 671.84 172.71 ;
   RECT 0.0 172.71 671.84 174.42 ;
   RECT 0.0 174.42 671.84 176.13 ;
   RECT 0.0 176.13 671.84 177.84 ;
   RECT 0.0 177.84 671.84 179.55 ;
   RECT 0.0 179.55 671.84 181.26 ;
   RECT 0.0 181.26 671.84 182.97 ;
   RECT 0.0 182.97 695.02 184.68 ;
   RECT 0.0 184.68 695.02 186.39 ;
   RECT 0.0 186.39 695.02 188.1 ;
   RECT 0.0 188.1 695.02 189.81 ;
   RECT 0.0 189.81 695.02 191.52 ;
   RECT 0.0 191.52 695.02 193.23 ;
   RECT 0.0 193.23 695.02 194.94 ;
   RECT 0.0 194.94 695.02 196.65 ;
   RECT 0.0 196.65 695.02 198.36 ;
   RECT 0.0 198.36 695.02 200.07 ;
   RECT 0.0 200.07 695.02 201.78 ;
   RECT 0.0 201.78 695.02 203.49 ;
   RECT 0.0 203.49 695.02 205.2 ;
   RECT 0.0 205.2 695.02 206.91 ;
   RECT 0.0 206.91 695.02 208.62 ;
   RECT 0.0 208.62 695.02 210.33 ;
   RECT 0.0 210.33 695.02 212.04 ;
   RECT 0.0 212.04 671.84 213.75 ;
   RECT 0.0 213.75 671.84 215.46 ;
   RECT 0.0 215.46 671.84 217.17 ;
   RECT 0.0 217.17 671.84 218.88 ;
   RECT 0.0 218.88 671.84 220.59 ;
   RECT 0.0 220.59 671.84 222.3 ;
   RECT 0.0 222.3 671.84 224.01 ;
   RECT 0.0 224.01 671.84 225.72 ;
   RECT 0.0 225.72 671.84 227.43 ;
   RECT 0.0 227.43 671.84 229.14 ;
   RECT 0.0 229.14 671.84 230.85 ;
   RECT 0.0 230.85 671.84 232.56 ;
   RECT 0.0 232.56 671.84 234.27 ;
   RECT 0.0 234.27 671.84 235.98 ;
   RECT 0.0 235.98 671.84 237.69 ;
   RECT 0.0 237.69 671.84 239.4 ;
   RECT 0.0 239.4 671.84 241.11 ;
   RECT 0.0 241.11 671.84 242.82 ;
   RECT 0.0 242.82 671.84 244.53 ;
   RECT 0.0 244.53 671.84 246.24 ;
   RECT 0.0 246.24 671.84 247.95 ;
   RECT 0.0 247.95 671.84 249.66 ;
   RECT 0.0 249.66 671.84 251.37 ;
   RECT 0.0 251.37 671.84 253.08 ;
   RECT 0.0 253.08 671.84 254.79 ;
   RECT 0.0 254.79 671.84 256.5 ;
   RECT 0.0 256.5 671.84 258.21 ;
   RECT 0.0 258.21 671.84 259.92 ;
   RECT 0.0 259.92 671.84 261.63 ;
   RECT 0.0 261.63 671.84 263.34 ;
   RECT 0.0 263.34 671.84 265.05 ;
   RECT 0.0 265.05 671.84 266.76 ;
   RECT 0.0 266.76 671.84 268.47 ;
   RECT 0.0 268.47 671.84 270.18 ;
   RECT 0.0 270.18 671.84 271.89 ;
   RECT 0.0 271.89 671.84 273.6 ;
   RECT 0.0 273.6 671.84 275.31 ;
   RECT 0.0 275.31 671.84 277.02 ;
   RECT 0.0 277.02 671.84 278.73 ;
   RECT 0.0 278.73 671.84 280.44 ;
   RECT 0.0 280.44 671.84 282.15 ;
   RECT 0.0 282.15 671.84 283.86 ;
   RECT 0.0 283.86 671.84 285.57 ;
   RECT 0.0 285.57 671.84 287.28 ;
   RECT 0.0 287.28 671.84 288.99 ;
   RECT 0.0 288.99 671.84 290.7 ;
   RECT 0.0 290.7 671.84 292.41 ;
   RECT 0.0 292.41 671.84 294.12 ;
   RECT 0.0 294.12 671.84 295.83 ;
   RECT 0.0 295.83 671.84 297.54 ;
   RECT 0.0 297.54 671.84 299.25 ;
   RECT 0.0 299.25 671.84 300.96 ;
   RECT 0.0 300.96 671.84 302.67 ;
   RECT 0.0 302.67 671.84 304.38 ;
   RECT 0.0 304.38 671.84 306.09 ;
   RECT 0.0 306.09 671.84 307.8 ;
   RECT 0.0 307.8 671.84 309.51 ;
   RECT 0.0 309.51 671.84 311.22 ;
   RECT 0.0 311.22 671.84 312.93 ;
   RECT 0.0 312.93 671.84 314.64 ;
   RECT 0.0 314.64 671.84 316.35 ;
   RECT 0.0 316.35 671.84 318.06 ;
   RECT 0.0 318.06 671.84 319.77 ;
   RECT 0.0 319.77 671.84 321.48 ;
   RECT 0.0 321.48 671.84 323.19 ;
   RECT 0.0 323.19 671.84 324.9 ;
   RECT 0.0 324.9 671.84 326.61 ;
   RECT 0.0 326.61 671.84 328.32 ;
   RECT 0.0 328.32 671.84 330.03 ;
   RECT 0.0 330.03 671.84 331.74 ;
   RECT 0.0 331.74 671.84 333.45 ;
   RECT 0.0 333.45 671.84 335.16 ;
   RECT 0.0 335.16 671.84 336.87 ;
   RECT 0.0 336.87 671.84 338.58 ;
   RECT 0.0 338.58 671.84 340.29 ;
   RECT 0.0 340.29 671.84 342.0 ;
   RECT 0.0 342.0 671.84 343.71 ;
   RECT 0.0 343.71 671.84 345.42 ;
   RECT 0.0 345.42 671.84 347.13 ;
   RECT 0.0 347.13 671.84 348.84 ;
   RECT 0.0 348.84 671.84 350.55 ;
   RECT 0.0 350.55 671.84 352.26 ;
   RECT 0.0 352.26 671.84 353.97 ;
   RECT 0.0 353.97 671.84 355.68 ;
   RECT 0.0 355.68 671.84 357.39 ;
   RECT 0.0 357.39 671.84 359.1 ;
   RECT 0.0 359.1 671.84 360.81 ;
   RECT 0.0 360.81 671.84 362.52 ;
   RECT 0.0 362.52 671.84 364.23 ;
   RECT 0.0 364.23 671.84 365.94 ;
   RECT 0.0 365.94 671.84 367.65 ;
   RECT 0.0 367.65 671.84 369.36 ;
   RECT 0.0 369.36 671.84 371.07 ;
   RECT 0.0 371.07 671.84 372.78 ;
   RECT 0.0 372.78 671.84 374.49 ;
   RECT 0.0 374.49 671.84 376.2 ;
   RECT 0.0 376.2 671.84 377.91 ;
   RECT 0.0 377.91 671.84 379.62 ;
   RECT 0.0 379.62 671.84 381.33 ;
   RECT 0.0 381.33 671.84 383.04 ;
   RECT 0.0 383.04 671.84 384.75 ;
   RECT 0.0 384.75 671.84 386.46 ;
   RECT 0.0 386.46 671.84 388.17 ;
   RECT 0.0 388.17 671.84 389.88 ;
   RECT 0.0 389.88 671.84 391.59 ;
   RECT 0.0 391.59 671.84 393.3 ;
   RECT 0.0 393.3 671.84 395.01 ;
   RECT 0.0 395.01 671.84 396.72 ;
   RECT 0.0 396.72 671.84 398.43 ;
   RECT 0.0 398.43 671.84 400.14 ;
   RECT 0.0 400.14 671.84 401.85 ;
   RECT 0.0 401.85 671.84 403.56 ;
   RECT 0.0 403.56 671.84 405.27 ;
   RECT 0.0 405.27 671.84 406.98 ;
   RECT 0.0 406.98 671.84 408.69 ;
   RECT 0.0 408.69 671.84 410.4 ;
  LAYER via1 ;
   RECT 0.0 0.0 671.84 1.71 ;
   RECT 0.0 1.71 671.84 3.42 ;
   RECT 0.0 3.42 671.84 5.13 ;
   RECT 0.0 5.13 671.84 6.84 ;
   RECT 0.0 6.84 671.84 8.55 ;
   RECT 0.0 8.55 671.84 10.26 ;
   RECT 0.0 10.26 671.84 11.97 ;
   RECT 0.0 11.97 671.84 13.68 ;
   RECT 0.0 13.68 671.84 15.39 ;
   RECT 0.0 15.39 671.84 17.1 ;
   RECT 0.0 17.1 671.84 18.81 ;
   RECT 0.0 18.81 671.84 20.52 ;
   RECT 0.0 20.52 671.84 22.23 ;
   RECT 0.0 22.23 671.84 23.94 ;
   RECT 0.0 23.94 671.84 25.65 ;
   RECT 0.0 25.65 671.84 27.36 ;
   RECT 0.0 27.36 671.84 29.07 ;
   RECT 0.0 29.07 671.84 30.78 ;
   RECT 0.0 30.78 671.84 32.49 ;
   RECT 0.0 32.49 671.84 34.2 ;
   RECT 0.0 34.2 671.84 35.91 ;
   RECT 0.0 35.91 671.84 37.62 ;
   RECT 0.0 37.62 671.84 39.33 ;
   RECT 0.0 39.33 671.84 41.04 ;
   RECT 0.0 41.04 671.84 42.75 ;
   RECT 0.0 42.75 671.84 44.46 ;
   RECT 0.0 44.46 671.84 46.17 ;
   RECT 0.0 46.17 671.84 47.88 ;
   RECT 0.0 47.88 671.84 49.59 ;
   RECT 0.0 49.59 671.84 51.3 ;
   RECT 0.0 51.3 671.84 53.01 ;
   RECT 0.0 53.01 671.84 54.72 ;
   RECT 0.0 54.72 671.84 56.43 ;
   RECT 0.0 56.43 671.84 58.14 ;
   RECT 0.0 58.14 671.84 59.85 ;
   RECT 0.0 59.85 671.84 61.56 ;
   RECT 0.0 61.56 671.84 63.27 ;
   RECT 0.0 63.27 671.84 64.98 ;
   RECT 0.0 64.98 671.84 66.69 ;
   RECT 0.0 66.69 671.84 68.4 ;
   RECT 0.0 68.4 671.84 70.11 ;
   RECT 0.0 70.11 671.84 71.82 ;
   RECT 0.0 71.82 671.84 73.53 ;
   RECT 0.0 73.53 671.84 75.24 ;
   RECT 0.0 75.24 671.84 76.95 ;
   RECT 0.0 76.95 671.84 78.66 ;
   RECT 0.0 78.66 671.84 80.37 ;
   RECT 0.0 80.37 671.84 82.08 ;
   RECT 0.0 82.08 671.84 83.79 ;
   RECT 0.0 83.79 671.84 85.5 ;
   RECT 0.0 85.5 671.84 87.21 ;
   RECT 0.0 87.21 671.84 88.92 ;
   RECT 0.0 88.92 671.84 90.63 ;
   RECT 0.0 90.63 671.84 92.34 ;
   RECT 0.0 92.34 671.84 94.05 ;
   RECT 0.0 94.05 671.84 95.76 ;
   RECT 0.0 95.76 671.84 97.47 ;
   RECT 0.0 97.47 671.84 99.18 ;
   RECT 0.0 99.18 671.84 100.89 ;
   RECT 0.0 100.89 671.84 102.6 ;
   RECT 0.0 102.6 671.84 104.31 ;
   RECT 0.0 104.31 671.84 106.02 ;
   RECT 0.0 106.02 671.84 107.73 ;
   RECT 0.0 107.73 671.84 109.44 ;
   RECT 0.0 109.44 671.84 111.15 ;
   RECT 0.0 111.15 671.84 112.86 ;
   RECT 0.0 112.86 671.84 114.57 ;
   RECT 0.0 114.57 671.84 116.28 ;
   RECT 0.0 116.28 671.84 117.99 ;
   RECT 0.0 117.99 671.84 119.7 ;
   RECT 0.0 119.7 671.84 121.41 ;
   RECT 0.0 121.41 671.84 123.12 ;
   RECT 0.0 123.12 671.84 124.83 ;
   RECT 0.0 124.83 671.84 126.54 ;
   RECT 0.0 126.54 671.84 128.25 ;
   RECT 0.0 128.25 671.84 129.96 ;
   RECT 0.0 129.96 671.84 131.67 ;
   RECT 0.0 131.67 671.84 133.38 ;
   RECT 0.0 133.38 671.84 135.09 ;
   RECT 0.0 135.09 671.84 136.8 ;
   RECT 0.0 136.8 671.84 138.51 ;
   RECT 0.0 138.51 671.84 140.22 ;
   RECT 0.0 140.22 671.84 141.93 ;
   RECT 0.0 141.93 671.84 143.64 ;
   RECT 0.0 143.64 671.84 145.35 ;
   RECT 0.0 145.35 671.84 147.06 ;
   RECT 0.0 147.06 671.84 148.77 ;
   RECT 0.0 148.77 671.84 150.48 ;
   RECT 0.0 150.48 671.84 152.19 ;
   RECT 0.0 152.19 671.84 153.9 ;
   RECT 0.0 153.9 671.84 155.61 ;
   RECT 0.0 155.61 671.84 157.32 ;
   RECT 0.0 157.32 671.84 159.03 ;
   RECT 0.0 159.03 671.84 160.74 ;
   RECT 0.0 160.74 671.84 162.45 ;
   RECT 0.0 162.45 671.84 164.16 ;
   RECT 0.0 164.16 671.84 165.87 ;
   RECT 0.0 165.87 671.84 167.58 ;
   RECT 0.0 167.58 671.84 169.29 ;
   RECT 0.0 169.29 671.84 171.0 ;
   RECT 0.0 171.0 671.84 172.71 ;
   RECT 0.0 172.71 671.84 174.42 ;
   RECT 0.0 174.42 671.84 176.13 ;
   RECT 0.0 176.13 671.84 177.84 ;
   RECT 0.0 177.84 671.84 179.55 ;
   RECT 0.0 179.55 671.84 181.26 ;
   RECT 0.0 181.26 671.84 182.97 ;
   RECT 0.0 182.97 695.02 184.68 ;
   RECT 0.0 184.68 695.02 186.39 ;
   RECT 0.0 186.39 695.02 188.1 ;
   RECT 0.0 188.1 695.02 189.81 ;
   RECT 0.0 189.81 695.02 191.52 ;
   RECT 0.0 191.52 695.02 193.23 ;
   RECT 0.0 193.23 695.02 194.94 ;
   RECT 0.0 194.94 695.02 196.65 ;
   RECT 0.0 196.65 695.02 198.36 ;
   RECT 0.0 198.36 695.02 200.07 ;
   RECT 0.0 200.07 695.02 201.78 ;
   RECT 0.0 201.78 695.02 203.49 ;
   RECT 0.0 203.49 695.02 205.2 ;
   RECT 0.0 205.2 695.02 206.91 ;
   RECT 0.0 206.91 695.02 208.62 ;
   RECT 0.0 208.62 695.02 210.33 ;
   RECT 0.0 210.33 695.02 212.04 ;
   RECT 0.0 212.04 671.84 213.75 ;
   RECT 0.0 213.75 671.84 215.46 ;
   RECT 0.0 215.46 671.84 217.17 ;
   RECT 0.0 217.17 671.84 218.88 ;
   RECT 0.0 218.88 671.84 220.59 ;
   RECT 0.0 220.59 671.84 222.3 ;
   RECT 0.0 222.3 671.84 224.01 ;
   RECT 0.0 224.01 671.84 225.72 ;
   RECT 0.0 225.72 671.84 227.43 ;
   RECT 0.0 227.43 671.84 229.14 ;
   RECT 0.0 229.14 671.84 230.85 ;
   RECT 0.0 230.85 671.84 232.56 ;
   RECT 0.0 232.56 671.84 234.27 ;
   RECT 0.0 234.27 671.84 235.98 ;
   RECT 0.0 235.98 671.84 237.69 ;
   RECT 0.0 237.69 671.84 239.4 ;
   RECT 0.0 239.4 671.84 241.11 ;
   RECT 0.0 241.11 671.84 242.82 ;
   RECT 0.0 242.82 671.84 244.53 ;
   RECT 0.0 244.53 671.84 246.24 ;
   RECT 0.0 246.24 671.84 247.95 ;
   RECT 0.0 247.95 671.84 249.66 ;
   RECT 0.0 249.66 671.84 251.37 ;
   RECT 0.0 251.37 671.84 253.08 ;
   RECT 0.0 253.08 671.84 254.79 ;
   RECT 0.0 254.79 671.84 256.5 ;
   RECT 0.0 256.5 671.84 258.21 ;
   RECT 0.0 258.21 671.84 259.92 ;
   RECT 0.0 259.92 671.84 261.63 ;
   RECT 0.0 261.63 671.84 263.34 ;
   RECT 0.0 263.34 671.84 265.05 ;
   RECT 0.0 265.05 671.84 266.76 ;
   RECT 0.0 266.76 671.84 268.47 ;
   RECT 0.0 268.47 671.84 270.18 ;
   RECT 0.0 270.18 671.84 271.89 ;
   RECT 0.0 271.89 671.84 273.6 ;
   RECT 0.0 273.6 671.84 275.31 ;
   RECT 0.0 275.31 671.84 277.02 ;
   RECT 0.0 277.02 671.84 278.73 ;
   RECT 0.0 278.73 671.84 280.44 ;
   RECT 0.0 280.44 671.84 282.15 ;
   RECT 0.0 282.15 671.84 283.86 ;
   RECT 0.0 283.86 671.84 285.57 ;
   RECT 0.0 285.57 671.84 287.28 ;
   RECT 0.0 287.28 671.84 288.99 ;
   RECT 0.0 288.99 671.84 290.7 ;
   RECT 0.0 290.7 671.84 292.41 ;
   RECT 0.0 292.41 671.84 294.12 ;
   RECT 0.0 294.12 671.84 295.83 ;
   RECT 0.0 295.83 671.84 297.54 ;
   RECT 0.0 297.54 671.84 299.25 ;
   RECT 0.0 299.25 671.84 300.96 ;
   RECT 0.0 300.96 671.84 302.67 ;
   RECT 0.0 302.67 671.84 304.38 ;
   RECT 0.0 304.38 671.84 306.09 ;
   RECT 0.0 306.09 671.84 307.8 ;
   RECT 0.0 307.8 671.84 309.51 ;
   RECT 0.0 309.51 671.84 311.22 ;
   RECT 0.0 311.22 671.84 312.93 ;
   RECT 0.0 312.93 671.84 314.64 ;
   RECT 0.0 314.64 671.84 316.35 ;
   RECT 0.0 316.35 671.84 318.06 ;
   RECT 0.0 318.06 671.84 319.77 ;
   RECT 0.0 319.77 671.84 321.48 ;
   RECT 0.0 321.48 671.84 323.19 ;
   RECT 0.0 323.19 671.84 324.9 ;
   RECT 0.0 324.9 671.84 326.61 ;
   RECT 0.0 326.61 671.84 328.32 ;
   RECT 0.0 328.32 671.84 330.03 ;
   RECT 0.0 330.03 671.84 331.74 ;
   RECT 0.0 331.74 671.84 333.45 ;
   RECT 0.0 333.45 671.84 335.16 ;
   RECT 0.0 335.16 671.84 336.87 ;
   RECT 0.0 336.87 671.84 338.58 ;
   RECT 0.0 338.58 671.84 340.29 ;
   RECT 0.0 340.29 671.84 342.0 ;
   RECT 0.0 342.0 671.84 343.71 ;
   RECT 0.0 343.71 671.84 345.42 ;
   RECT 0.0 345.42 671.84 347.13 ;
   RECT 0.0 347.13 671.84 348.84 ;
   RECT 0.0 348.84 671.84 350.55 ;
   RECT 0.0 350.55 671.84 352.26 ;
   RECT 0.0 352.26 671.84 353.97 ;
   RECT 0.0 353.97 671.84 355.68 ;
   RECT 0.0 355.68 671.84 357.39 ;
   RECT 0.0 357.39 671.84 359.1 ;
   RECT 0.0 359.1 671.84 360.81 ;
   RECT 0.0 360.81 671.84 362.52 ;
   RECT 0.0 362.52 671.84 364.23 ;
   RECT 0.0 364.23 671.84 365.94 ;
   RECT 0.0 365.94 671.84 367.65 ;
   RECT 0.0 367.65 671.84 369.36 ;
   RECT 0.0 369.36 671.84 371.07 ;
   RECT 0.0 371.07 671.84 372.78 ;
   RECT 0.0 372.78 671.84 374.49 ;
   RECT 0.0 374.49 671.84 376.2 ;
   RECT 0.0 376.2 671.84 377.91 ;
   RECT 0.0 377.91 671.84 379.62 ;
   RECT 0.0 379.62 671.84 381.33 ;
   RECT 0.0 381.33 671.84 383.04 ;
   RECT 0.0 383.04 671.84 384.75 ;
   RECT 0.0 384.75 671.84 386.46 ;
   RECT 0.0 386.46 671.84 388.17 ;
   RECT 0.0 388.17 671.84 389.88 ;
   RECT 0.0 389.88 671.84 391.59 ;
   RECT 0.0 391.59 671.84 393.3 ;
   RECT 0.0 393.3 671.84 395.01 ;
   RECT 0.0 395.01 671.84 396.72 ;
   RECT 0.0 396.72 671.84 398.43 ;
   RECT 0.0 398.43 671.84 400.14 ;
   RECT 0.0 400.14 671.84 401.85 ;
   RECT 0.0 401.85 671.84 403.56 ;
   RECT 0.0 403.56 671.84 405.27 ;
   RECT 0.0 405.27 671.84 406.98 ;
   RECT 0.0 406.98 671.84 408.69 ;
   RECT 0.0 408.69 671.84 410.4 ;
  LAYER metal2 ;
   RECT 0.0 0.0 671.84 1.71 ;
   RECT 0.0 1.71 671.84 3.42 ;
   RECT 0.0 3.42 671.84 5.13 ;
   RECT 0.0 5.13 671.84 6.84 ;
   RECT 0.0 6.84 671.84 8.55 ;
   RECT 0.0 8.55 671.84 10.26 ;
   RECT 0.0 10.26 671.84 11.97 ;
   RECT 0.0 11.97 671.84 13.68 ;
   RECT 0.0 13.68 671.84 15.39 ;
   RECT 0.0 15.39 671.84 17.1 ;
   RECT 0.0 17.1 671.84 18.81 ;
   RECT 0.0 18.81 671.84 20.52 ;
   RECT 0.0 20.52 671.84 22.23 ;
   RECT 0.0 22.23 671.84 23.94 ;
   RECT 0.0 23.94 671.84 25.65 ;
   RECT 0.0 25.65 671.84 27.36 ;
   RECT 0.0 27.36 671.84 29.07 ;
   RECT 0.0 29.07 671.84 30.78 ;
   RECT 0.0 30.78 671.84 32.49 ;
   RECT 0.0 32.49 671.84 34.2 ;
   RECT 0.0 34.2 671.84 35.91 ;
   RECT 0.0 35.91 671.84 37.62 ;
   RECT 0.0 37.62 671.84 39.33 ;
   RECT 0.0 39.33 671.84 41.04 ;
   RECT 0.0 41.04 671.84 42.75 ;
   RECT 0.0 42.75 671.84 44.46 ;
   RECT 0.0 44.46 671.84 46.17 ;
   RECT 0.0 46.17 671.84 47.88 ;
   RECT 0.0 47.88 671.84 49.59 ;
   RECT 0.0 49.59 671.84 51.3 ;
   RECT 0.0 51.3 671.84 53.01 ;
   RECT 0.0 53.01 671.84 54.72 ;
   RECT 0.0 54.72 671.84 56.43 ;
   RECT 0.0 56.43 671.84 58.14 ;
   RECT 0.0 58.14 671.84 59.85 ;
   RECT 0.0 59.85 671.84 61.56 ;
   RECT 0.0 61.56 671.84 63.27 ;
   RECT 0.0 63.27 671.84 64.98 ;
   RECT 0.0 64.98 671.84 66.69 ;
   RECT 0.0 66.69 671.84 68.4 ;
   RECT 0.0 68.4 671.84 70.11 ;
   RECT 0.0 70.11 671.84 71.82 ;
   RECT 0.0 71.82 671.84 73.53 ;
   RECT 0.0 73.53 671.84 75.24 ;
   RECT 0.0 75.24 671.84 76.95 ;
   RECT 0.0 76.95 671.84 78.66 ;
   RECT 0.0 78.66 671.84 80.37 ;
   RECT 0.0 80.37 671.84 82.08 ;
   RECT 0.0 82.08 671.84 83.79 ;
   RECT 0.0 83.79 671.84 85.5 ;
   RECT 0.0 85.5 671.84 87.21 ;
   RECT 0.0 87.21 671.84 88.92 ;
   RECT 0.0 88.92 671.84 90.63 ;
   RECT 0.0 90.63 671.84 92.34 ;
   RECT 0.0 92.34 671.84 94.05 ;
   RECT 0.0 94.05 671.84 95.76 ;
   RECT 0.0 95.76 671.84 97.47 ;
   RECT 0.0 97.47 671.84 99.18 ;
   RECT 0.0 99.18 671.84 100.89 ;
   RECT 0.0 100.89 671.84 102.6 ;
   RECT 0.0 102.6 671.84 104.31 ;
   RECT 0.0 104.31 671.84 106.02 ;
   RECT 0.0 106.02 671.84 107.73 ;
   RECT 0.0 107.73 671.84 109.44 ;
   RECT 0.0 109.44 671.84 111.15 ;
   RECT 0.0 111.15 671.84 112.86 ;
   RECT 0.0 112.86 671.84 114.57 ;
   RECT 0.0 114.57 671.84 116.28 ;
   RECT 0.0 116.28 671.84 117.99 ;
   RECT 0.0 117.99 671.84 119.7 ;
   RECT 0.0 119.7 671.84 121.41 ;
   RECT 0.0 121.41 671.84 123.12 ;
   RECT 0.0 123.12 671.84 124.83 ;
   RECT 0.0 124.83 671.84 126.54 ;
   RECT 0.0 126.54 671.84 128.25 ;
   RECT 0.0 128.25 671.84 129.96 ;
   RECT 0.0 129.96 671.84 131.67 ;
   RECT 0.0 131.67 671.84 133.38 ;
   RECT 0.0 133.38 671.84 135.09 ;
   RECT 0.0 135.09 671.84 136.8 ;
   RECT 0.0 136.8 671.84 138.51 ;
   RECT 0.0 138.51 671.84 140.22 ;
   RECT 0.0 140.22 671.84 141.93 ;
   RECT 0.0 141.93 671.84 143.64 ;
   RECT 0.0 143.64 671.84 145.35 ;
   RECT 0.0 145.35 671.84 147.06 ;
   RECT 0.0 147.06 671.84 148.77 ;
   RECT 0.0 148.77 671.84 150.48 ;
   RECT 0.0 150.48 671.84 152.19 ;
   RECT 0.0 152.19 671.84 153.9 ;
   RECT 0.0 153.9 671.84 155.61 ;
   RECT 0.0 155.61 671.84 157.32 ;
   RECT 0.0 157.32 671.84 159.03 ;
   RECT 0.0 159.03 671.84 160.74 ;
   RECT 0.0 160.74 671.84 162.45 ;
   RECT 0.0 162.45 671.84 164.16 ;
   RECT 0.0 164.16 671.84 165.87 ;
   RECT 0.0 165.87 671.84 167.58 ;
   RECT 0.0 167.58 671.84 169.29 ;
   RECT 0.0 169.29 671.84 171.0 ;
   RECT 0.0 171.0 671.84 172.71 ;
   RECT 0.0 172.71 671.84 174.42 ;
   RECT 0.0 174.42 671.84 176.13 ;
   RECT 0.0 176.13 671.84 177.84 ;
   RECT 0.0 177.84 671.84 179.55 ;
   RECT 0.0 179.55 671.84 181.26 ;
   RECT 0.0 181.26 671.84 182.97 ;
   RECT 0.0 182.97 695.02 184.68 ;
   RECT 0.0 184.68 695.02 186.39 ;
   RECT 0.0 186.39 695.02 188.1 ;
   RECT 0.0 188.1 695.02 189.81 ;
   RECT 0.0 189.81 695.02 191.52 ;
   RECT 0.0 191.52 695.02 193.23 ;
   RECT 0.0 193.23 695.02 194.94 ;
   RECT 0.0 194.94 695.02 196.65 ;
   RECT 0.0 196.65 695.02 198.36 ;
   RECT 0.0 198.36 695.02 200.07 ;
   RECT 0.0 200.07 695.02 201.78 ;
   RECT 0.0 201.78 695.02 203.49 ;
   RECT 0.0 203.49 695.02 205.2 ;
   RECT 0.0 205.2 695.02 206.91 ;
   RECT 0.0 206.91 695.02 208.62 ;
   RECT 0.0 208.62 695.02 210.33 ;
   RECT 0.0 210.33 695.02 212.04 ;
   RECT 0.0 212.04 671.84 213.75 ;
   RECT 0.0 213.75 671.84 215.46 ;
   RECT 0.0 215.46 671.84 217.17 ;
   RECT 0.0 217.17 671.84 218.88 ;
   RECT 0.0 218.88 671.84 220.59 ;
   RECT 0.0 220.59 671.84 222.3 ;
   RECT 0.0 222.3 671.84 224.01 ;
   RECT 0.0 224.01 671.84 225.72 ;
   RECT 0.0 225.72 671.84 227.43 ;
   RECT 0.0 227.43 671.84 229.14 ;
   RECT 0.0 229.14 671.84 230.85 ;
   RECT 0.0 230.85 671.84 232.56 ;
   RECT 0.0 232.56 671.84 234.27 ;
   RECT 0.0 234.27 671.84 235.98 ;
   RECT 0.0 235.98 671.84 237.69 ;
   RECT 0.0 237.69 671.84 239.4 ;
   RECT 0.0 239.4 671.84 241.11 ;
   RECT 0.0 241.11 671.84 242.82 ;
   RECT 0.0 242.82 671.84 244.53 ;
   RECT 0.0 244.53 671.84 246.24 ;
   RECT 0.0 246.24 671.84 247.95 ;
   RECT 0.0 247.95 671.84 249.66 ;
   RECT 0.0 249.66 671.84 251.37 ;
   RECT 0.0 251.37 671.84 253.08 ;
   RECT 0.0 253.08 671.84 254.79 ;
   RECT 0.0 254.79 671.84 256.5 ;
   RECT 0.0 256.5 671.84 258.21 ;
   RECT 0.0 258.21 671.84 259.92 ;
   RECT 0.0 259.92 671.84 261.63 ;
   RECT 0.0 261.63 671.84 263.34 ;
   RECT 0.0 263.34 671.84 265.05 ;
   RECT 0.0 265.05 671.84 266.76 ;
   RECT 0.0 266.76 671.84 268.47 ;
   RECT 0.0 268.47 671.84 270.18 ;
   RECT 0.0 270.18 671.84 271.89 ;
   RECT 0.0 271.89 671.84 273.6 ;
   RECT 0.0 273.6 671.84 275.31 ;
   RECT 0.0 275.31 671.84 277.02 ;
   RECT 0.0 277.02 671.84 278.73 ;
   RECT 0.0 278.73 671.84 280.44 ;
   RECT 0.0 280.44 671.84 282.15 ;
   RECT 0.0 282.15 671.84 283.86 ;
   RECT 0.0 283.86 671.84 285.57 ;
   RECT 0.0 285.57 671.84 287.28 ;
   RECT 0.0 287.28 671.84 288.99 ;
   RECT 0.0 288.99 671.84 290.7 ;
   RECT 0.0 290.7 671.84 292.41 ;
   RECT 0.0 292.41 671.84 294.12 ;
   RECT 0.0 294.12 671.84 295.83 ;
   RECT 0.0 295.83 671.84 297.54 ;
   RECT 0.0 297.54 671.84 299.25 ;
   RECT 0.0 299.25 671.84 300.96 ;
   RECT 0.0 300.96 671.84 302.67 ;
   RECT 0.0 302.67 671.84 304.38 ;
   RECT 0.0 304.38 671.84 306.09 ;
   RECT 0.0 306.09 671.84 307.8 ;
   RECT 0.0 307.8 671.84 309.51 ;
   RECT 0.0 309.51 671.84 311.22 ;
   RECT 0.0 311.22 671.84 312.93 ;
   RECT 0.0 312.93 671.84 314.64 ;
   RECT 0.0 314.64 671.84 316.35 ;
   RECT 0.0 316.35 671.84 318.06 ;
   RECT 0.0 318.06 671.84 319.77 ;
   RECT 0.0 319.77 671.84 321.48 ;
   RECT 0.0 321.48 671.84 323.19 ;
   RECT 0.0 323.19 671.84 324.9 ;
   RECT 0.0 324.9 671.84 326.61 ;
   RECT 0.0 326.61 671.84 328.32 ;
   RECT 0.0 328.32 671.84 330.03 ;
   RECT 0.0 330.03 671.84 331.74 ;
   RECT 0.0 331.74 671.84 333.45 ;
   RECT 0.0 333.45 671.84 335.16 ;
   RECT 0.0 335.16 671.84 336.87 ;
   RECT 0.0 336.87 671.84 338.58 ;
   RECT 0.0 338.58 671.84 340.29 ;
   RECT 0.0 340.29 671.84 342.0 ;
   RECT 0.0 342.0 671.84 343.71 ;
   RECT 0.0 343.71 671.84 345.42 ;
   RECT 0.0 345.42 671.84 347.13 ;
   RECT 0.0 347.13 671.84 348.84 ;
   RECT 0.0 348.84 671.84 350.55 ;
   RECT 0.0 350.55 671.84 352.26 ;
   RECT 0.0 352.26 671.84 353.97 ;
   RECT 0.0 353.97 671.84 355.68 ;
   RECT 0.0 355.68 671.84 357.39 ;
   RECT 0.0 357.39 671.84 359.1 ;
   RECT 0.0 359.1 671.84 360.81 ;
   RECT 0.0 360.81 671.84 362.52 ;
   RECT 0.0 362.52 671.84 364.23 ;
   RECT 0.0 364.23 671.84 365.94 ;
   RECT 0.0 365.94 671.84 367.65 ;
   RECT 0.0 367.65 671.84 369.36 ;
   RECT 0.0 369.36 671.84 371.07 ;
   RECT 0.0 371.07 671.84 372.78 ;
   RECT 0.0 372.78 671.84 374.49 ;
   RECT 0.0 374.49 671.84 376.2 ;
   RECT 0.0 376.2 671.84 377.91 ;
   RECT 0.0 377.91 671.84 379.62 ;
   RECT 0.0 379.62 671.84 381.33 ;
   RECT 0.0 381.33 671.84 383.04 ;
   RECT 0.0 383.04 671.84 384.75 ;
   RECT 0.0 384.75 671.84 386.46 ;
   RECT 0.0 386.46 671.84 388.17 ;
   RECT 0.0 388.17 671.84 389.88 ;
   RECT 0.0 389.88 671.84 391.59 ;
   RECT 0.0 391.59 671.84 393.3 ;
   RECT 0.0 393.3 671.84 395.01 ;
   RECT 0.0 395.01 671.84 396.72 ;
   RECT 0.0 396.72 671.84 398.43 ;
   RECT 0.0 398.43 671.84 400.14 ;
   RECT 0.0 400.14 671.84 401.85 ;
   RECT 0.0 401.85 671.84 403.56 ;
   RECT 0.0 403.56 671.84 405.27 ;
   RECT 0.0 405.27 671.84 406.98 ;
   RECT 0.0 406.98 671.84 408.69 ;
   RECT 0.0 408.69 671.84 410.4 ;
  LAYER via2 ;
   RECT 0.0 0.0 671.84 1.71 ;
   RECT 0.0 1.71 671.84 3.42 ;
   RECT 0.0 3.42 671.84 5.13 ;
   RECT 0.0 5.13 671.84 6.84 ;
   RECT 0.0 6.84 671.84 8.55 ;
   RECT 0.0 8.55 671.84 10.26 ;
   RECT 0.0 10.26 671.84 11.97 ;
   RECT 0.0 11.97 671.84 13.68 ;
   RECT 0.0 13.68 671.84 15.39 ;
   RECT 0.0 15.39 671.84 17.1 ;
   RECT 0.0 17.1 671.84 18.81 ;
   RECT 0.0 18.81 671.84 20.52 ;
   RECT 0.0 20.52 671.84 22.23 ;
   RECT 0.0 22.23 671.84 23.94 ;
   RECT 0.0 23.94 671.84 25.65 ;
   RECT 0.0 25.65 671.84 27.36 ;
   RECT 0.0 27.36 671.84 29.07 ;
   RECT 0.0 29.07 671.84 30.78 ;
   RECT 0.0 30.78 671.84 32.49 ;
   RECT 0.0 32.49 671.84 34.2 ;
   RECT 0.0 34.2 671.84 35.91 ;
   RECT 0.0 35.91 671.84 37.62 ;
   RECT 0.0 37.62 671.84 39.33 ;
   RECT 0.0 39.33 671.84 41.04 ;
   RECT 0.0 41.04 671.84 42.75 ;
   RECT 0.0 42.75 671.84 44.46 ;
   RECT 0.0 44.46 671.84 46.17 ;
   RECT 0.0 46.17 671.84 47.88 ;
   RECT 0.0 47.88 671.84 49.59 ;
   RECT 0.0 49.59 671.84 51.3 ;
   RECT 0.0 51.3 671.84 53.01 ;
   RECT 0.0 53.01 671.84 54.72 ;
   RECT 0.0 54.72 671.84 56.43 ;
   RECT 0.0 56.43 671.84 58.14 ;
   RECT 0.0 58.14 671.84 59.85 ;
   RECT 0.0 59.85 671.84 61.56 ;
   RECT 0.0 61.56 671.84 63.27 ;
   RECT 0.0 63.27 671.84 64.98 ;
   RECT 0.0 64.98 671.84 66.69 ;
   RECT 0.0 66.69 671.84 68.4 ;
   RECT 0.0 68.4 671.84 70.11 ;
   RECT 0.0 70.11 671.84 71.82 ;
   RECT 0.0 71.82 671.84 73.53 ;
   RECT 0.0 73.53 671.84 75.24 ;
   RECT 0.0 75.24 671.84 76.95 ;
   RECT 0.0 76.95 671.84 78.66 ;
   RECT 0.0 78.66 671.84 80.37 ;
   RECT 0.0 80.37 671.84 82.08 ;
   RECT 0.0 82.08 671.84 83.79 ;
   RECT 0.0 83.79 671.84 85.5 ;
   RECT 0.0 85.5 671.84 87.21 ;
   RECT 0.0 87.21 671.84 88.92 ;
   RECT 0.0 88.92 671.84 90.63 ;
   RECT 0.0 90.63 671.84 92.34 ;
   RECT 0.0 92.34 671.84 94.05 ;
   RECT 0.0 94.05 671.84 95.76 ;
   RECT 0.0 95.76 671.84 97.47 ;
   RECT 0.0 97.47 671.84 99.18 ;
   RECT 0.0 99.18 671.84 100.89 ;
   RECT 0.0 100.89 671.84 102.6 ;
   RECT 0.0 102.6 671.84 104.31 ;
   RECT 0.0 104.31 671.84 106.02 ;
   RECT 0.0 106.02 671.84 107.73 ;
   RECT 0.0 107.73 671.84 109.44 ;
   RECT 0.0 109.44 671.84 111.15 ;
   RECT 0.0 111.15 671.84 112.86 ;
   RECT 0.0 112.86 671.84 114.57 ;
   RECT 0.0 114.57 671.84 116.28 ;
   RECT 0.0 116.28 671.84 117.99 ;
   RECT 0.0 117.99 671.84 119.7 ;
   RECT 0.0 119.7 671.84 121.41 ;
   RECT 0.0 121.41 671.84 123.12 ;
   RECT 0.0 123.12 671.84 124.83 ;
   RECT 0.0 124.83 671.84 126.54 ;
   RECT 0.0 126.54 671.84 128.25 ;
   RECT 0.0 128.25 671.84 129.96 ;
   RECT 0.0 129.96 671.84 131.67 ;
   RECT 0.0 131.67 671.84 133.38 ;
   RECT 0.0 133.38 671.84 135.09 ;
   RECT 0.0 135.09 671.84 136.8 ;
   RECT 0.0 136.8 671.84 138.51 ;
   RECT 0.0 138.51 671.84 140.22 ;
   RECT 0.0 140.22 671.84 141.93 ;
   RECT 0.0 141.93 671.84 143.64 ;
   RECT 0.0 143.64 671.84 145.35 ;
   RECT 0.0 145.35 671.84 147.06 ;
   RECT 0.0 147.06 671.84 148.77 ;
   RECT 0.0 148.77 671.84 150.48 ;
   RECT 0.0 150.48 671.84 152.19 ;
   RECT 0.0 152.19 671.84 153.9 ;
   RECT 0.0 153.9 671.84 155.61 ;
   RECT 0.0 155.61 671.84 157.32 ;
   RECT 0.0 157.32 671.84 159.03 ;
   RECT 0.0 159.03 671.84 160.74 ;
   RECT 0.0 160.74 671.84 162.45 ;
   RECT 0.0 162.45 671.84 164.16 ;
   RECT 0.0 164.16 671.84 165.87 ;
   RECT 0.0 165.87 671.84 167.58 ;
   RECT 0.0 167.58 671.84 169.29 ;
   RECT 0.0 169.29 671.84 171.0 ;
   RECT 0.0 171.0 671.84 172.71 ;
   RECT 0.0 172.71 671.84 174.42 ;
   RECT 0.0 174.42 671.84 176.13 ;
   RECT 0.0 176.13 671.84 177.84 ;
   RECT 0.0 177.84 671.84 179.55 ;
   RECT 0.0 179.55 671.84 181.26 ;
   RECT 0.0 181.26 671.84 182.97 ;
   RECT 0.0 182.97 695.02 184.68 ;
   RECT 0.0 184.68 695.02 186.39 ;
   RECT 0.0 186.39 695.02 188.1 ;
   RECT 0.0 188.1 695.02 189.81 ;
   RECT 0.0 189.81 695.02 191.52 ;
   RECT 0.0 191.52 695.02 193.23 ;
   RECT 0.0 193.23 695.02 194.94 ;
   RECT 0.0 194.94 695.02 196.65 ;
   RECT 0.0 196.65 695.02 198.36 ;
   RECT 0.0 198.36 695.02 200.07 ;
   RECT 0.0 200.07 695.02 201.78 ;
   RECT 0.0 201.78 695.02 203.49 ;
   RECT 0.0 203.49 695.02 205.2 ;
   RECT 0.0 205.2 695.02 206.91 ;
   RECT 0.0 206.91 695.02 208.62 ;
   RECT 0.0 208.62 695.02 210.33 ;
   RECT 0.0 210.33 695.02 212.04 ;
   RECT 0.0 212.04 671.84 213.75 ;
   RECT 0.0 213.75 671.84 215.46 ;
   RECT 0.0 215.46 671.84 217.17 ;
   RECT 0.0 217.17 671.84 218.88 ;
   RECT 0.0 218.88 671.84 220.59 ;
   RECT 0.0 220.59 671.84 222.3 ;
   RECT 0.0 222.3 671.84 224.01 ;
   RECT 0.0 224.01 671.84 225.72 ;
   RECT 0.0 225.72 671.84 227.43 ;
   RECT 0.0 227.43 671.84 229.14 ;
   RECT 0.0 229.14 671.84 230.85 ;
   RECT 0.0 230.85 671.84 232.56 ;
   RECT 0.0 232.56 671.84 234.27 ;
   RECT 0.0 234.27 671.84 235.98 ;
   RECT 0.0 235.98 671.84 237.69 ;
   RECT 0.0 237.69 671.84 239.4 ;
   RECT 0.0 239.4 671.84 241.11 ;
   RECT 0.0 241.11 671.84 242.82 ;
   RECT 0.0 242.82 671.84 244.53 ;
   RECT 0.0 244.53 671.84 246.24 ;
   RECT 0.0 246.24 671.84 247.95 ;
   RECT 0.0 247.95 671.84 249.66 ;
   RECT 0.0 249.66 671.84 251.37 ;
   RECT 0.0 251.37 671.84 253.08 ;
   RECT 0.0 253.08 671.84 254.79 ;
   RECT 0.0 254.79 671.84 256.5 ;
   RECT 0.0 256.5 671.84 258.21 ;
   RECT 0.0 258.21 671.84 259.92 ;
   RECT 0.0 259.92 671.84 261.63 ;
   RECT 0.0 261.63 671.84 263.34 ;
   RECT 0.0 263.34 671.84 265.05 ;
   RECT 0.0 265.05 671.84 266.76 ;
   RECT 0.0 266.76 671.84 268.47 ;
   RECT 0.0 268.47 671.84 270.18 ;
   RECT 0.0 270.18 671.84 271.89 ;
   RECT 0.0 271.89 671.84 273.6 ;
   RECT 0.0 273.6 671.84 275.31 ;
   RECT 0.0 275.31 671.84 277.02 ;
   RECT 0.0 277.02 671.84 278.73 ;
   RECT 0.0 278.73 671.84 280.44 ;
   RECT 0.0 280.44 671.84 282.15 ;
   RECT 0.0 282.15 671.84 283.86 ;
   RECT 0.0 283.86 671.84 285.57 ;
   RECT 0.0 285.57 671.84 287.28 ;
   RECT 0.0 287.28 671.84 288.99 ;
   RECT 0.0 288.99 671.84 290.7 ;
   RECT 0.0 290.7 671.84 292.41 ;
   RECT 0.0 292.41 671.84 294.12 ;
   RECT 0.0 294.12 671.84 295.83 ;
   RECT 0.0 295.83 671.84 297.54 ;
   RECT 0.0 297.54 671.84 299.25 ;
   RECT 0.0 299.25 671.84 300.96 ;
   RECT 0.0 300.96 671.84 302.67 ;
   RECT 0.0 302.67 671.84 304.38 ;
   RECT 0.0 304.38 671.84 306.09 ;
   RECT 0.0 306.09 671.84 307.8 ;
   RECT 0.0 307.8 671.84 309.51 ;
   RECT 0.0 309.51 671.84 311.22 ;
   RECT 0.0 311.22 671.84 312.93 ;
   RECT 0.0 312.93 671.84 314.64 ;
   RECT 0.0 314.64 671.84 316.35 ;
   RECT 0.0 316.35 671.84 318.06 ;
   RECT 0.0 318.06 671.84 319.77 ;
   RECT 0.0 319.77 671.84 321.48 ;
   RECT 0.0 321.48 671.84 323.19 ;
   RECT 0.0 323.19 671.84 324.9 ;
   RECT 0.0 324.9 671.84 326.61 ;
   RECT 0.0 326.61 671.84 328.32 ;
   RECT 0.0 328.32 671.84 330.03 ;
   RECT 0.0 330.03 671.84 331.74 ;
   RECT 0.0 331.74 671.84 333.45 ;
   RECT 0.0 333.45 671.84 335.16 ;
   RECT 0.0 335.16 671.84 336.87 ;
   RECT 0.0 336.87 671.84 338.58 ;
   RECT 0.0 338.58 671.84 340.29 ;
   RECT 0.0 340.29 671.84 342.0 ;
   RECT 0.0 342.0 671.84 343.71 ;
   RECT 0.0 343.71 671.84 345.42 ;
   RECT 0.0 345.42 671.84 347.13 ;
   RECT 0.0 347.13 671.84 348.84 ;
   RECT 0.0 348.84 671.84 350.55 ;
   RECT 0.0 350.55 671.84 352.26 ;
   RECT 0.0 352.26 671.84 353.97 ;
   RECT 0.0 353.97 671.84 355.68 ;
   RECT 0.0 355.68 671.84 357.39 ;
   RECT 0.0 357.39 671.84 359.1 ;
   RECT 0.0 359.1 671.84 360.81 ;
   RECT 0.0 360.81 671.84 362.52 ;
   RECT 0.0 362.52 671.84 364.23 ;
   RECT 0.0 364.23 671.84 365.94 ;
   RECT 0.0 365.94 671.84 367.65 ;
   RECT 0.0 367.65 671.84 369.36 ;
   RECT 0.0 369.36 671.84 371.07 ;
   RECT 0.0 371.07 671.84 372.78 ;
   RECT 0.0 372.78 671.84 374.49 ;
   RECT 0.0 374.49 671.84 376.2 ;
   RECT 0.0 376.2 671.84 377.91 ;
   RECT 0.0 377.91 671.84 379.62 ;
   RECT 0.0 379.62 671.84 381.33 ;
   RECT 0.0 381.33 671.84 383.04 ;
   RECT 0.0 383.04 671.84 384.75 ;
   RECT 0.0 384.75 671.84 386.46 ;
   RECT 0.0 386.46 671.84 388.17 ;
   RECT 0.0 388.17 671.84 389.88 ;
   RECT 0.0 389.88 671.84 391.59 ;
   RECT 0.0 391.59 671.84 393.3 ;
   RECT 0.0 393.3 671.84 395.01 ;
   RECT 0.0 395.01 671.84 396.72 ;
   RECT 0.0 396.72 671.84 398.43 ;
   RECT 0.0 398.43 671.84 400.14 ;
   RECT 0.0 400.14 671.84 401.85 ;
   RECT 0.0 401.85 671.84 403.56 ;
   RECT 0.0 403.56 671.84 405.27 ;
   RECT 0.0 405.27 671.84 406.98 ;
   RECT 0.0 406.98 671.84 408.69 ;
   RECT 0.0 408.69 671.84 410.4 ;
  LAYER metal3 ;
   RECT 0.0 0.0 671.84 1.71 ;
   RECT 0.0 1.71 671.84 3.42 ;
   RECT 0.0 3.42 671.84 5.13 ;
   RECT 0.0 5.13 671.84 6.84 ;
   RECT 0.0 6.84 671.84 8.55 ;
   RECT 0.0 8.55 671.84 10.26 ;
   RECT 0.0 10.26 671.84 11.97 ;
   RECT 0.0 11.97 671.84 13.68 ;
   RECT 0.0 13.68 671.84 15.39 ;
   RECT 0.0 15.39 671.84 17.1 ;
   RECT 0.0 17.1 671.84 18.81 ;
   RECT 0.0 18.81 671.84 20.52 ;
   RECT 0.0 20.52 671.84 22.23 ;
   RECT 0.0 22.23 671.84 23.94 ;
   RECT 0.0 23.94 671.84 25.65 ;
   RECT 0.0 25.65 671.84 27.36 ;
   RECT 0.0 27.36 671.84 29.07 ;
   RECT 0.0 29.07 671.84 30.78 ;
   RECT 0.0 30.78 671.84 32.49 ;
   RECT 0.0 32.49 671.84 34.2 ;
   RECT 0.0 34.2 671.84 35.91 ;
   RECT 0.0 35.91 671.84 37.62 ;
   RECT 0.0 37.62 671.84 39.33 ;
   RECT 0.0 39.33 671.84 41.04 ;
   RECT 0.0 41.04 671.84 42.75 ;
   RECT 0.0 42.75 671.84 44.46 ;
   RECT 0.0 44.46 671.84 46.17 ;
   RECT 0.0 46.17 671.84 47.88 ;
   RECT 0.0 47.88 671.84 49.59 ;
   RECT 0.0 49.59 671.84 51.3 ;
   RECT 0.0 51.3 671.84 53.01 ;
   RECT 0.0 53.01 671.84 54.72 ;
   RECT 0.0 54.72 671.84 56.43 ;
   RECT 0.0 56.43 671.84 58.14 ;
   RECT 0.0 58.14 671.84 59.85 ;
   RECT 0.0 59.85 671.84 61.56 ;
   RECT 0.0 61.56 671.84 63.27 ;
   RECT 0.0 63.27 671.84 64.98 ;
   RECT 0.0 64.98 671.84 66.69 ;
   RECT 0.0 66.69 671.84 68.4 ;
   RECT 0.0 68.4 671.84 70.11 ;
   RECT 0.0 70.11 671.84 71.82 ;
   RECT 0.0 71.82 671.84 73.53 ;
   RECT 0.0 73.53 671.84 75.24 ;
   RECT 0.0 75.24 671.84 76.95 ;
   RECT 0.0 76.95 671.84 78.66 ;
   RECT 0.0 78.66 671.84 80.37 ;
   RECT 0.0 80.37 671.84 82.08 ;
   RECT 0.0 82.08 671.84 83.79 ;
   RECT 0.0 83.79 671.84 85.5 ;
   RECT 0.0 85.5 671.84 87.21 ;
   RECT 0.0 87.21 671.84 88.92 ;
   RECT 0.0 88.92 671.84 90.63 ;
   RECT 0.0 90.63 671.84 92.34 ;
   RECT 0.0 92.34 671.84 94.05 ;
   RECT 0.0 94.05 671.84 95.76 ;
   RECT 0.0 95.76 671.84 97.47 ;
   RECT 0.0 97.47 671.84 99.18 ;
   RECT 0.0 99.18 671.84 100.89 ;
   RECT 0.0 100.89 671.84 102.6 ;
   RECT 0.0 102.6 671.84 104.31 ;
   RECT 0.0 104.31 671.84 106.02 ;
   RECT 0.0 106.02 671.84 107.73 ;
   RECT 0.0 107.73 671.84 109.44 ;
   RECT 0.0 109.44 671.84 111.15 ;
   RECT 0.0 111.15 671.84 112.86 ;
   RECT 0.0 112.86 671.84 114.57 ;
   RECT 0.0 114.57 671.84 116.28 ;
   RECT 0.0 116.28 671.84 117.99 ;
   RECT 0.0 117.99 671.84 119.7 ;
   RECT 0.0 119.7 671.84 121.41 ;
   RECT 0.0 121.41 671.84 123.12 ;
   RECT 0.0 123.12 671.84 124.83 ;
   RECT 0.0 124.83 671.84 126.54 ;
   RECT 0.0 126.54 671.84 128.25 ;
   RECT 0.0 128.25 671.84 129.96 ;
   RECT 0.0 129.96 671.84 131.67 ;
   RECT 0.0 131.67 671.84 133.38 ;
   RECT 0.0 133.38 671.84 135.09 ;
   RECT 0.0 135.09 671.84 136.8 ;
   RECT 0.0 136.8 671.84 138.51 ;
   RECT 0.0 138.51 671.84 140.22 ;
   RECT 0.0 140.22 671.84 141.93 ;
   RECT 0.0 141.93 671.84 143.64 ;
   RECT 0.0 143.64 671.84 145.35 ;
   RECT 0.0 145.35 671.84 147.06 ;
   RECT 0.0 147.06 671.84 148.77 ;
   RECT 0.0 148.77 671.84 150.48 ;
   RECT 0.0 150.48 671.84 152.19 ;
   RECT 0.0 152.19 671.84 153.9 ;
   RECT 0.0 153.9 671.84 155.61 ;
   RECT 0.0 155.61 671.84 157.32 ;
   RECT 0.0 157.32 671.84 159.03 ;
   RECT 0.0 159.03 671.84 160.74 ;
   RECT 0.0 160.74 671.84 162.45 ;
   RECT 0.0 162.45 671.84 164.16 ;
   RECT 0.0 164.16 671.84 165.87 ;
   RECT 0.0 165.87 671.84 167.58 ;
   RECT 0.0 167.58 671.84 169.29 ;
   RECT 0.0 169.29 671.84 171.0 ;
   RECT 0.0 171.0 671.84 172.71 ;
   RECT 0.0 172.71 671.84 174.42 ;
   RECT 0.0 174.42 671.84 176.13 ;
   RECT 0.0 176.13 671.84 177.84 ;
   RECT 0.0 177.84 671.84 179.55 ;
   RECT 0.0 179.55 671.84 181.26 ;
   RECT 0.0 181.26 671.84 182.97 ;
   RECT 0.0 182.97 695.02 184.68 ;
   RECT 0.0 184.68 695.02 186.39 ;
   RECT 0.0 186.39 695.02 188.1 ;
   RECT 0.0 188.1 695.02 189.81 ;
   RECT 0.0 189.81 695.02 191.52 ;
   RECT 0.0 191.52 695.02 193.23 ;
   RECT 0.0 193.23 695.02 194.94 ;
   RECT 0.0 194.94 695.02 196.65 ;
   RECT 0.0 196.65 695.02 198.36 ;
   RECT 0.0 198.36 695.02 200.07 ;
   RECT 0.0 200.07 695.02 201.78 ;
   RECT 0.0 201.78 695.02 203.49 ;
   RECT 0.0 203.49 695.02 205.2 ;
   RECT 0.0 205.2 695.02 206.91 ;
   RECT 0.0 206.91 695.02 208.62 ;
   RECT 0.0 208.62 695.02 210.33 ;
   RECT 0.0 210.33 695.02 212.04 ;
   RECT 0.0 212.04 671.84 213.75 ;
   RECT 0.0 213.75 671.84 215.46 ;
   RECT 0.0 215.46 671.84 217.17 ;
   RECT 0.0 217.17 671.84 218.88 ;
   RECT 0.0 218.88 671.84 220.59 ;
   RECT 0.0 220.59 671.84 222.3 ;
   RECT 0.0 222.3 671.84 224.01 ;
   RECT 0.0 224.01 671.84 225.72 ;
   RECT 0.0 225.72 671.84 227.43 ;
   RECT 0.0 227.43 671.84 229.14 ;
   RECT 0.0 229.14 671.84 230.85 ;
   RECT 0.0 230.85 671.84 232.56 ;
   RECT 0.0 232.56 671.84 234.27 ;
   RECT 0.0 234.27 671.84 235.98 ;
   RECT 0.0 235.98 671.84 237.69 ;
   RECT 0.0 237.69 671.84 239.4 ;
   RECT 0.0 239.4 671.84 241.11 ;
   RECT 0.0 241.11 671.84 242.82 ;
   RECT 0.0 242.82 671.84 244.53 ;
   RECT 0.0 244.53 671.84 246.24 ;
   RECT 0.0 246.24 671.84 247.95 ;
   RECT 0.0 247.95 671.84 249.66 ;
   RECT 0.0 249.66 671.84 251.37 ;
   RECT 0.0 251.37 671.84 253.08 ;
   RECT 0.0 253.08 671.84 254.79 ;
   RECT 0.0 254.79 671.84 256.5 ;
   RECT 0.0 256.5 671.84 258.21 ;
   RECT 0.0 258.21 671.84 259.92 ;
   RECT 0.0 259.92 671.84 261.63 ;
   RECT 0.0 261.63 671.84 263.34 ;
   RECT 0.0 263.34 671.84 265.05 ;
   RECT 0.0 265.05 671.84 266.76 ;
   RECT 0.0 266.76 671.84 268.47 ;
   RECT 0.0 268.47 671.84 270.18 ;
   RECT 0.0 270.18 671.84 271.89 ;
   RECT 0.0 271.89 671.84 273.6 ;
   RECT 0.0 273.6 671.84 275.31 ;
   RECT 0.0 275.31 671.84 277.02 ;
   RECT 0.0 277.02 671.84 278.73 ;
   RECT 0.0 278.73 671.84 280.44 ;
   RECT 0.0 280.44 671.84 282.15 ;
   RECT 0.0 282.15 671.84 283.86 ;
   RECT 0.0 283.86 671.84 285.57 ;
   RECT 0.0 285.57 671.84 287.28 ;
   RECT 0.0 287.28 671.84 288.99 ;
   RECT 0.0 288.99 671.84 290.7 ;
   RECT 0.0 290.7 671.84 292.41 ;
   RECT 0.0 292.41 671.84 294.12 ;
   RECT 0.0 294.12 671.84 295.83 ;
   RECT 0.0 295.83 671.84 297.54 ;
   RECT 0.0 297.54 671.84 299.25 ;
   RECT 0.0 299.25 671.84 300.96 ;
   RECT 0.0 300.96 671.84 302.67 ;
   RECT 0.0 302.67 671.84 304.38 ;
   RECT 0.0 304.38 671.84 306.09 ;
   RECT 0.0 306.09 671.84 307.8 ;
   RECT 0.0 307.8 671.84 309.51 ;
   RECT 0.0 309.51 671.84 311.22 ;
   RECT 0.0 311.22 671.84 312.93 ;
   RECT 0.0 312.93 671.84 314.64 ;
   RECT 0.0 314.64 671.84 316.35 ;
   RECT 0.0 316.35 671.84 318.06 ;
   RECT 0.0 318.06 671.84 319.77 ;
   RECT 0.0 319.77 671.84 321.48 ;
   RECT 0.0 321.48 671.84 323.19 ;
   RECT 0.0 323.19 671.84 324.9 ;
   RECT 0.0 324.9 671.84 326.61 ;
   RECT 0.0 326.61 671.84 328.32 ;
   RECT 0.0 328.32 671.84 330.03 ;
   RECT 0.0 330.03 671.84 331.74 ;
   RECT 0.0 331.74 671.84 333.45 ;
   RECT 0.0 333.45 671.84 335.16 ;
   RECT 0.0 335.16 671.84 336.87 ;
   RECT 0.0 336.87 671.84 338.58 ;
   RECT 0.0 338.58 671.84 340.29 ;
   RECT 0.0 340.29 671.84 342.0 ;
   RECT 0.0 342.0 671.84 343.71 ;
   RECT 0.0 343.71 671.84 345.42 ;
   RECT 0.0 345.42 671.84 347.13 ;
   RECT 0.0 347.13 671.84 348.84 ;
   RECT 0.0 348.84 671.84 350.55 ;
   RECT 0.0 350.55 671.84 352.26 ;
   RECT 0.0 352.26 671.84 353.97 ;
   RECT 0.0 353.97 671.84 355.68 ;
   RECT 0.0 355.68 671.84 357.39 ;
   RECT 0.0 357.39 671.84 359.1 ;
   RECT 0.0 359.1 671.84 360.81 ;
   RECT 0.0 360.81 671.84 362.52 ;
   RECT 0.0 362.52 671.84 364.23 ;
   RECT 0.0 364.23 671.84 365.94 ;
   RECT 0.0 365.94 671.84 367.65 ;
   RECT 0.0 367.65 671.84 369.36 ;
   RECT 0.0 369.36 671.84 371.07 ;
   RECT 0.0 371.07 671.84 372.78 ;
   RECT 0.0 372.78 671.84 374.49 ;
   RECT 0.0 374.49 671.84 376.2 ;
   RECT 0.0 376.2 671.84 377.91 ;
   RECT 0.0 377.91 671.84 379.62 ;
   RECT 0.0 379.62 671.84 381.33 ;
   RECT 0.0 381.33 671.84 383.04 ;
   RECT 0.0 383.04 671.84 384.75 ;
   RECT 0.0 384.75 671.84 386.46 ;
   RECT 0.0 386.46 671.84 388.17 ;
   RECT 0.0 388.17 671.84 389.88 ;
   RECT 0.0 389.88 671.84 391.59 ;
   RECT 0.0 391.59 671.84 393.3 ;
   RECT 0.0 393.3 671.84 395.01 ;
   RECT 0.0 395.01 671.84 396.72 ;
   RECT 0.0 396.72 671.84 398.43 ;
   RECT 0.0 398.43 671.84 400.14 ;
   RECT 0.0 400.14 671.84 401.85 ;
   RECT 0.0 401.85 671.84 403.56 ;
   RECT 0.0 403.56 671.84 405.27 ;
   RECT 0.0 405.27 671.84 406.98 ;
   RECT 0.0 406.98 671.84 408.69 ;
   RECT 0.0 408.69 671.84 410.4 ;
  LAYER via3 ;
   RECT 0.0 0.0 671.84 1.71 ;
   RECT 0.0 1.71 671.84 3.42 ;
   RECT 0.0 3.42 671.84 5.13 ;
   RECT 0.0 5.13 671.84 6.84 ;
   RECT 0.0 6.84 671.84 8.55 ;
   RECT 0.0 8.55 671.84 10.26 ;
   RECT 0.0 10.26 671.84 11.97 ;
   RECT 0.0 11.97 671.84 13.68 ;
   RECT 0.0 13.68 671.84 15.39 ;
   RECT 0.0 15.39 671.84 17.1 ;
   RECT 0.0 17.1 671.84 18.81 ;
   RECT 0.0 18.81 671.84 20.52 ;
   RECT 0.0 20.52 671.84 22.23 ;
   RECT 0.0 22.23 671.84 23.94 ;
   RECT 0.0 23.94 671.84 25.65 ;
   RECT 0.0 25.65 671.84 27.36 ;
   RECT 0.0 27.36 671.84 29.07 ;
   RECT 0.0 29.07 671.84 30.78 ;
   RECT 0.0 30.78 671.84 32.49 ;
   RECT 0.0 32.49 671.84 34.2 ;
   RECT 0.0 34.2 671.84 35.91 ;
   RECT 0.0 35.91 671.84 37.62 ;
   RECT 0.0 37.62 671.84 39.33 ;
   RECT 0.0 39.33 671.84 41.04 ;
   RECT 0.0 41.04 671.84 42.75 ;
   RECT 0.0 42.75 671.84 44.46 ;
   RECT 0.0 44.46 671.84 46.17 ;
   RECT 0.0 46.17 671.84 47.88 ;
   RECT 0.0 47.88 671.84 49.59 ;
   RECT 0.0 49.59 671.84 51.3 ;
   RECT 0.0 51.3 671.84 53.01 ;
   RECT 0.0 53.01 671.84 54.72 ;
   RECT 0.0 54.72 671.84 56.43 ;
   RECT 0.0 56.43 671.84 58.14 ;
   RECT 0.0 58.14 671.84 59.85 ;
   RECT 0.0 59.85 671.84 61.56 ;
   RECT 0.0 61.56 671.84 63.27 ;
   RECT 0.0 63.27 671.84 64.98 ;
   RECT 0.0 64.98 671.84 66.69 ;
   RECT 0.0 66.69 671.84 68.4 ;
   RECT 0.0 68.4 671.84 70.11 ;
   RECT 0.0 70.11 671.84 71.82 ;
   RECT 0.0 71.82 671.84 73.53 ;
   RECT 0.0 73.53 671.84 75.24 ;
   RECT 0.0 75.24 671.84 76.95 ;
   RECT 0.0 76.95 671.84 78.66 ;
   RECT 0.0 78.66 671.84 80.37 ;
   RECT 0.0 80.37 671.84 82.08 ;
   RECT 0.0 82.08 671.84 83.79 ;
   RECT 0.0 83.79 671.84 85.5 ;
   RECT 0.0 85.5 671.84 87.21 ;
   RECT 0.0 87.21 671.84 88.92 ;
   RECT 0.0 88.92 671.84 90.63 ;
   RECT 0.0 90.63 671.84 92.34 ;
   RECT 0.0 92.34 671.84 94.05 ;
   RECT 0.0 94.05 671.84 95.76 ;
   RECT 0.0 95.76 671.84 97.47 ;
   RECT 0.0 97.47 671.84 99.18 ;
   RECT 0.0 99.18 671.84 100.89 ;
   RECT 0.0 100.89 671.84 102.6 ;
   RECT 0.0 102.6 671.84 104.31 ;
   RECT 0.0 104.31 671.84 106.02 ;
   RECT 0.0 106.02 671.84 107.73 ;
   RECT 0.0 107.73 671.84 109.44 ;
   RECT 0.0 109.44 671.84 111.15 ;
   RECT 0.0 111.15 671.84 112.86 ;
   RECT 0.0 112.86 671.84 114.57 ;
   RECT 0.0 114.57 671.84 116.28 ;
   RECT 0.0 116.28 671.84 117.99 ;
   RECT 0.0 117.99 671.84 119.7 ;
   RECT 0.0 119.7 671.84 121.41 ;
   RECT 0.0 121.41 671.84 123.12 ;
   RECT 0.0 123.12 671.84 124.83 ;
   RECT 0.0 124.83 671.84 126.54 ;
   RECT 0.0 126.54 671.84 128.25 ;
   RECT 0.0 128.25 671.84 129.96 ;
   RECT 0.0 129.96 671.84 131.67 ;
   RECT 0.0 131.67 671.84 133.38 ;
   RECT 0.0 133.38 671.84 135.09 ;
   RECT 0.0 135.09 671.84 136.8 ;
   RECT 0.0 136.8 671.84 138.51 ;
   RECT 0.0 138.51 671.84 140.22 ;
   RECT 0.0 140.22 671.84 141.93 ;
   RECT 0.0 141.93 671.84 143.64 ;
   RECT 0.0 143.64 671.84 145.35 ;
   RECT 0.0 145.35 671.84 147.06 ;
   RECT 0.0 147.06 671.84 148.77 ;
   RECT 0.0 148.77 671.84 150.48 ;
   RECT 0.0 150.48 671.84 152.19 ;
   RECT 0.0 152.19 671.84 153.9 ;
   RECT 0.0 153.9 671.84 155.61 ;
   RECT 0.0 155.61 671.84 157.32 ;
   RECT 0.0 157.32 671.84 159.03 ;
   RECT 0.0 159.03 671.84 160.74 ;
   RECT 0.0 160.74 671.84 162.45 ;
   RECT 0.0 162.45 671.84 164.16 ;
   RECT 0.0 164.16 671.84 165.87 ;
   RECT 0.0 165.87 671.84 167.58 ;
   RECT 0.0 167.58 671.84 169.29 ;
   RECT 0.0 169.29 671.84 171.0 ;
   RECT 0.0 171.0 671.84 172.71 ;
   RECT 0.0 172.71 671.84 174.42 ;
   RECT 0.0 174.42 671.84 176.13 ;
   RECT 0.0 176.13 671.84 177.84 ;
   RECT 0.0 177.84 671.84 179.55 ;
   RECT 0.0 179.55 671.84 181.26 ;
   RECT 0.0 181.26 671.84 182.97 ;
   RECT 0.0 182.97 695.02 184.68 ;
   RECT 0.0 184.68 695.02 186.39 ;
   RECT 0.0 186.39 695.02 188.1 ;
   RECT 0.0 188.1 695.02 189.81 ;
   RECT 0.0 189.81 695.02 191.52 ;
   RECT 0.0 191.52 695.02 193.23 ;
   RECT 0.0 193.23 695.02 194.94 ;
   RECT 0.0 194.94 695.02 196.65 ;
   RECT 0.0 196.65 695.02 198.36 ;
   RECT 0.0 198.36 695.02 200.07 ;
   RECT 0.0 200.07 695.02 201.78 ;
   RECT 0.0 201.78 695.02 203.49 ;
   RECT 0.0 203.49 695.02 205.2 ;
   RECT 0.0 205.2 695.02 206.91 ;
   RECT 0.0 206.91 695.02 208.62 ;
   RECT 0.0 208.62 695.02 210.33 ;
   RECT 0.0 210.33 695.02 212.04 ;
   RECT 0.0 212.04 671.84 213.75 ;
   RECT 0.0 213.75 671.84 215.46 ;
   RECT 0.0 215.46 671.84 217.17 ;
   RECT 0.0 217.17 671.84 218.88 ;
   RECT 0.0 218.88 671.84 220.59 ;
   RECT 0.0 220.59 671.84 222.3 ;
   RECT 0.0 222.3 671.84 224.01 ;
   RECT 0.0 224.01 671.84 225.72 ;
   RECT 0.0 225.72 671.84 227.43 ;
   RECT 0.0 227.43 671.84 229.14 ;
   RECT 0.0 229.14 671.84 230.85 ;
   RECT 0.0 230.85 671.84 232.56 ;
   RECT 0.0 232.56 671.84 234.27 ;
   RECT 0.0 234.27 671.84 235.98 ;
   RECT 0.0 235.98 671.84 237.69 ;
   RECT 0.0 237.69 671.84 239.4 ;
   RECT 0.0 239.4 671.84 241.11 ;
   RECT 0.0 241.11 671.84 242.82 ;
   RECT 0.0 242.82 671.84 244.53 ;
   RECT 0.0 244.53 671.84 246.24 ;
   RECT 0.0 246.24 671.84 247.95 ;
   RECT 0.0 247.95 671.84 249.66 ;
   RECT 0.0 249.66 671.84 251.37 ;
   RECT 0.0 251.37 671.84 253.08 ;
   RECT 0.0 253.08 671.84 254.79 ;
   RECT 0.0 254.79 671.84 256.5 ;
   RECT 0.0 256.5 671.84 258.21 ;
   RECT 0.0 258.21 671.84 259.92 ;
   RECT 0.0 259.92 671.84 261.63 ;
   RECT 0.0 261.63 671.84 263.34 ;
   RECT 0.0 263.34 671.84 265.05 ;
   RECT 0.0 265.05 671.84 266.76 ;
   RECT 0.0 266.76 671.84 268.47 ;
   RECT 0.0 268.47 671.84 270.18 ;
   RECT 0.0 270.18 671.84 271.89 ;
   RECT 0.0 271.89 671.84 273.6 ;
   RECT 0.0 273.6 671.84 275.31 ;
   RECT 0.0 275.31 671.84 277.02 ;
   RECT 0.0 277.02 671.84 278.73 ;
   RECT 0.0 278.73 671.84 280.44 ;
   RECT 0.0 280.44 671.84 282.15 ;
   RECT 0.0 282.15 671.84 283.86 ;
   RECT 0.0 283.86 671.84 285.57 ;
   RECT 0.0 285.57 671.84 287.28 ;
   RECT 0.0 287.28 671.84 288.99 ;
   RECT 0.0 288.99 671.84 290.7 ;
   RECT 0.0 290.7 671.84 292.41 ;
   RECT 0.0 292.41 671.84 294.12 ;
   RECT 0.0 294.12 671.84 295.83 ;
   RECT 0.0 295.83 671.84 297.54 ;
   RECT 0.0 297.54 671.84 299.25 ;
   RECT 0.0 299.25 671.84 300.96 ;
   RECT 0.0 300.96 671.84 302.67 ;
   RECT 0.0 302.67 671.84 304.38 ;
   RECT 0.0 304.38 671.84 306.09 ;
   RECT 0.0 306.09 671.84 307.8 ;
   RECT 0.0 307.8 671.84 309.51 ;
   RECT 0.0 309.51 671.84 311.22 ;
   RECT 0.0 311.22 671.84 312.93 ;
   RECT 0.0 312.93 671.84 314.64 ;
   RECT 0.0 314.64 671.84 316.35 ;
   RECT 0.0 316.35 671.84 318.06 ;
   RECT 0.0 318.06 671.84 319.77 ;
   RECT 0.0 319.77 671.84 321.48 ;
   RECT 0.0 321.48 671.84 323.19 ;
   RECT 0.0 323.19 671.84 324.9 ;
   RECT 0.0 324.9 671.84 326.61 ;
   RECT 0.0 326.61 671.84 328.32 ;
   RECT 0.0 328.32 671.84 330.03 ;
   RECT 0.0 330.03 671.84 331.74 ;
   RECT 0.0 331.74 671.84 333.45 ;
   RECT 0.0 333.45 671.84 335.16 ;
   RECT 0.0 335.16 671.84 336.87 ;
   RECT 0.0 336.87 671.84 338.58 ;
   RECT 0.0 338.58 671.84 340.29 ;
   RECT 0.0 340.29 671.84 342.0 ;
   RECT 0.0 342.0 671.84 343.71 ;
   RECT 0.0 343.71 671.84 345.42 ;
   RECT 0.0 345.42 671.84 347.13 ;
   RECT 0.0 347.13 671.84 348.84 ;
   RECT 0.0 348.84 671.84 350.55 ;
   RECT 0.0 350.55 671.84 352.26 ;
   RECT 0.0 352.26 671.84 353.97 ;
   RECT 0.0 353.97 671.84 355.68 ;
   RECT 0.0 355.68 671.84 357.39 ;
   RECT 0.0 357.39 671.84 359.1 ;
   RECT 0.0 359.1 671.84 360.81 ;
   RECT 0.0 360.81 671.84 362.52 ;
   RECT 0.0 362.52 671.84 364.23 ;
   RECT 0.0 364.23 671.84 365.94 ;
   RECT 0.0 365.94 671.84 367.65 ;
   RECT 0.0 367.65 671.84 369.36 ;
   RECT 0.0 369.36 671.84 371.07 ;
   RECT 0.0 371.07 671.84 372.78 ;
   RECT 0.0 372.78 671.84 374.49 ;
   RECT 0.0 374.49 671.84 376.2 ;
   RECT 0.0 376.2 671.84 377.91 ;
   RECT 0.0 377.91 671.84 379.62 ;
   RECT 0.0 379.62 671.84 381.33 ;
   RECT 0.0 381.33 671.84 383.04 ;
   RECT 0.0 383.04 671.84 384.75 ;
   RECT 0.0 384.75 671.84 386.46 ;
   RECT 0.0 386.46 671.84 388.17 ;
   RECT 0.0 388.17 671.84 389.88 ;
   RECT 0.0 389.88 671.84 391.59 ;
   RECT 0.0 391.59 671.84 393.3 ;
   RECT 0.0 393.3 671.84 395.01 ;
   RECT 0.0 395.01 671.84 396.72 ;
   RECT 0.0 396.72 671.84 398.43 ;
   RECT 0.0 398.43 671.84 400.14 ;
   RECT 0.0 400.14 671.84 401.85 ;
   RECT 0.0 401.85 671.84 403.56 ;
   RECT 0.0 403.56 671.84 405.27 ;
   RECT 0.0 405.27 671.84 406.98 ;
   RECT 0.0 406.98 671.84 408.69 ;
   RECT 0.0 408.69 671.84 410.4 ;
  LAYER metal4 ;
   RECT 0.0 0.0 671.84 1.71 ;
   RECT 0.0 1.71 671.84 3.42 ;
   RECT 0.0 3.42 671.84 5.13 ;
   RECT 0.0 5.13 671.84 6.84 ;
   RECT 0.0 6.84 671.84 8.55 ;
   RECT 0.0 8.55 671.84 10.26 ;
   RECT 0.0 10.26 671.84 11.97 ;
   RECT 0.0 11.97 671.84 13.68 ;
   RECT 0.0 13.68 671.84 15.39 ;
   RECT 0.0 15.39 671.84 17.1 ;
   RECT 0.0 17.1 671.84 18.81 ;
   RECT 0.0 18.81 671.84 20.52 ;
   RECT 0.0 20.52 671.84 22.23 ;
   RECT 0.0 22.23 671.84 23.94 ;
   RECT 0.0 23.94 671.84 25.65 ;
   RECT 0.0 25.65 671.84 27.36 ;
   RECT 0.0 27.36 671.84 29.07 ;
   RECT 0.0 29.07 671.84 30.78 ;
   RECT 0.0 30.78 671.84 32.49 ;
   RECT 0.0 32.49 671.84 34.2 ;
   RECT 0.0 34.2 671.84 35.91 ;
   RECT 0.0 35.91 671.84 37.62 ;
   RECT 0.0 37.62 671.84 39.33 ;
   RECT 0.0 39.33 671.84 41.04 ;
   RECT 0.0 41.04 671.84 42.75 ;
   RECT 0.0 42.75 671.84 44.46 ;
   RECT 0.0 44.46 671.84 46.17 ;
   RECT 0.0 46.17 671.84 47.88 ;
   RECT 0.0 47.88 671.84 49.59 ;
   RECT 0.0 49.59 671.84 51.3 ;
   RECT 0.0 51.3 671.84 53.01 ;
   RECT 0.0 53.01 671.84 54.72 ;
   RECT 0.0 54.72 671.84 56.43 ;
   RECT 0.0 56.43 671.84 58.14 ;
   RECT 0.0 58.14 671.84 59.85 ;
   RECT 0.0 59.85 671.84 61.56 ;
   RECT 0.0 61.56 671.84 63.27 ;
   RECT 0.0 63.27 671.84 64.98 ;
   RECT 0.0 64.98 671.84 66.69 ;
   RECT 0.0 66.69 671.84 68.4 ;
   RECT 0.0 68.4 671.84 70.11 ;
   RECT 0.0 70.11 671.84 71.82 ;
   RECT 0.0 71.82 671.84 73.53 ;
   RECT 0.0 73.53 671.84 75.24 ;
   RECT 0.0 75.24 671.84 76.95 ;
   RECT 0.0 76.95 671.84 78.66 ;
   RECT 0.0 78.66 671.84 80.37 ;
   RECT 0.0 80.37 671.84 82.08 ;
   RECT 0.0 82.08 671.84 83.79 ;
   RECT 0.0 83.79 671.84 85.5 ;
   RECT 0.0 85.5 671.84 87.21 ;
   RECT 0.0 87.21 671.84 88.92 ;
   RECT 0.0 88.92 671.84 90.63 ;
   RECT 0.0 90.63 671.84 92.34 ;
   RECT 0.0 92.34 671.84 94.05 ;
   RECT 0.0 94.05 671.84 95.76 ;
   RECT 0.0 95.76 671.84 97.47 ;
   RECT 0.0 97.47 671.84 99.18 ;
   RECT 0.0 99.18 671.84 100.89 ;
   RECT 0.0 100.89 671.84 102.6 ;
   RECT 0.0 102.6 671.84 104.31 ;
   RECT 0.0 104.31 671.84 106.02 ;
   RECT 0.0 106.02 671.84 107.73 ;
   RECT 0.0 107.73 671.84 109.44 ;
   RECT 0.0 109.44 671.84 111.15 ;
   RECT 0.0 111.15 671.84 112.86 ;
   RECT 0.0 112.86 671.84 114.57 ;
   RECT 0.0 114.57 671.84 116.28 ;
   RECT 0.0 116.28 671.84 117.99 ;
   RECT 0.0 117.99 671.84 119.7 ;
   RECT 0.0 119.7 671.84 121.41 ;
   RECT 0.0 121.41 671.84 123.12 ;
   RECT 0.0 123.12 671.84 124.83 ;
   RECT 0.0 124.83 671.84 126.54 ;
   RECT 0.0 126.54 671.84 128.25 ;
   RECT 0.0 128.25 671.84 129.96 ;
   RECT 0.0 129.96 671.84 131.67 ;
   RECT 0.0 131.67 671.84 133.38 ;
   RECT 0.0 133.38 671.84 135.09 ;
   RECT 0.0 135.09 671.84 136.8 ;
   RECT 0.0 136.8 671.84 138.51 ;
   RECT 0.0 138.51 671.84 140.22 ;
   RECT 0.0 140.22 671.84 141.93 ;
   RECT 0.0 141.93 671.84 143.64 ;
   RECT 0.0 143.64 671.84 145.35 ;
   RECT 0.0 145.35 671.84 147.06 ;
   RECT 0.0 147.06 671.84 148.77 ;
   RECT 0.0 148.77 671.84 150.48 ;
   RECT 0.0 150.48 671.84 152.19 ;
   RECT 0.0 152.19 671.84 153.9 ;
   RECT 0.0 153.9 671.84 155.61 ;
   RECT 0.0 155.61 671.84 157.32 ;
   RECT 0.0 157.32 671.84 159.03 ;
   RECT 0.0 159.03 671.84 160.74 ;
   RECT 0.0 160.74 671.84 162.45 ;
   RECT 0.0 162.45 671.84 164.16 ;
   RECT 0.0 164.16 671.84 165.87 ;
   RECT 0.0 165.87 671.84 167.58 ;
   RECT 0.0 167.58 671.84 169.29 ;
   RECT 0.0 169.29 671.84 171.0 ;
   RECT 0.0 171.0 671.84 172.71 ;
   RECT 0.0 172.71 671.84 174.42 ;
   RECT 0.0 174.42 671.84 176.13 ;
   RECT 0.0 176.13 671.84 177.84 ;
   RECT 0.0 177.84 671.84 179.55 ;
   RECT 0.0 179.55 671.84 181.26 ;
   RECT 0.0 181.26 671.84 182.97 ;
   RECT 0.0 182.97 695.02 184.68 ;
   RECT 0.0 184.68 695.02 186.39 ;
   RECT 0.0 186.39 695.02 188.1 ;
   RECT 0.0 188.1 695.02 189.81 ;
   RECT 0.0 189.81 695.02 191.52 ;
   RECT 0.0 191.52 695.02 193.23 ;
   RECT 0.0 193.23 695.02 194.94 ;
   RECT 0.0 194.94 695.02 196.65 ;
   RECT 0.0 196.65 695.02 198.36 ;
   RECT 0.0 198.36 695.02 200.07 ;
   RECT 0.0 200.07 695.02 201.78 ;
   RECT 0.0 201.78 695.02 203.49 ;
   RECT 0.0 203.49 695.02 205.2 ;
   RECT 0.0 205.2 695.02 206.91 ;
   RECT 0.0 206.91 695.02 208.62 ;
   RECT 0.0 208.62 695.02 210.33 ;
   RECT 0.0 210.33 695.02 212.04 ;
   RECT 0.0 212.04 671.84 213.75 ;
   RECT 0.0 213.75 671.84 215.46 ;
   RECT 0.0 215.46 671.84 217.17 ;
   RECT 0.0 217.17 671.84 218.88 ;
   RECT 0.0 218.88 671.84 220.59 ;
   RECT 0.0 220.59 671.84 222.3 ;
   RECT 0.0 222.3 671.84 224.01 ;
   RECT 0.0 224.01 671.84 225.72 ;
   RECT 0.0 225.72 671.84 227.43 ;
   RECT 0.0 227.43 671.84 229.14 ;
   RECT 0.0 229.14 671.84 230.85 ;
   RECT 0.0 230.85 671.84 232.56 ;
   RECT 0.0 232.56 671.84 234.27 ;
   RECT 0.0 234.27 671.84 235.98 ;
   RECT 0.0 235.98 671.84 237.69 ;
   RECT 0.0 237.69 671.84 239.4 ;
   RECT 0.0 239.4 671.84 241.11 ;
   RECT 0.0 241.11 671.84 242.82 ;
   RECT 0.0 242.82 671.84 244.53 ;
   RECT 0.0 244.53 671.84 246.24 ;
   RECT 0.0 246.24 671.84 247.95 ;
   RECT 0.0 247.95 671.84 249.66 ;
   RECT 0.0 249.66 671.84 251.37 ;
   RECT 0.0 251.37 671.84 253.08 ;
   RECT 0.0 253.08 671.84 254.79 ;
   RECT 0.0 254.79 671.84 256.5 ;
   RECT 0.0 256.5 671.84 258.21 ;
   RECT 0.0 258.21 671.84 259.92 ;
   RECT 0.0 259.92 671.84 261.63 ;
   RECT 0.0 261.63 671.84 263.34 ;
   RECT 0.0 263.34 671.84 265.05 ;
   RECT 0.0 265.05 671.84 266.76 ;
   RECT 0.0 266.76 671.84 268.47 ;
   RECT 0.0 268.47 671.84 270.18 ;
   RECT 0.0 270.18 671.84 271.89 ;
   RECT 0.0 271.89 671.84 273.6 ;
   RECT 0.0 273.6 671.84 275.31 ;
   RECT 0.0 275.31 671.84 277.02 ;
   RECT 0.0 277.02 671.84 278.73 ;
   RECT 0.0 278.73 671.84 280.44 ;
   RECT 0.0 280.44 671.84 282.15 ;
   RECT 0.0 282.15 671.84 283.86 ;
   RECT 0.0 283.86 671.84 285.57 ;
   RECT 0.0 285.57 671.84 287.28 ;
   RECT 0.0 287.28 671.84 288.99 ;
   RECT 0.0 288.99 671.84 290.7 ;
   RECT 0.0 290.7 671.84 292.41 ;
   RECT 0.0 292.41 671.84 294.12 ;
   RECT 0.0 294.12 671.84 295.83 ;
   RECT 0.0 295.83 671.84 297.54 ;
   RECT 0.0 297.54 671.84 299.25 ;
   RECT 0.0 299.25 671.84 300.96 ;
   RECT 0.0 300.96 671.84 302.67 ;
   RECT 0.0 302.67 671.84 304.38 ;
   RECT 0.0 304.38 671.84 306.09 ;
   RECT 0.0 306.09 671.84 307.8 ;
   RECT 0.0 307.8 671.84 309.51 ;
   RECT 0.0 309.51 671.84 311.22 ;
   RECT 0.0 311.22 671.84 312.93 ;
   RECT 0.0 312.93 671.84 314.64 ;
   RECT 0.0 314.64 671.84 316.35 ;
   RECT 0.0 316.35 671.84 318.06 ;
   RECT 0.0 318.06 671.84 319.77 ;
   RECT 0.0 319.77 671.84 321.48 ;
   RECT 0.0 321.48 671.84 323.19 ;
   RECT 0.0 323.19 671.84 324.9 ;
   RECT 0.0 324.9 671.84 326.61 ;
   RECT 0.0 326.61 671.84 328.32 ;
   RECT 0.0 328.32 671.84 330.03 ;
   RECT 0.0 330.03 671.84 331.74 ;
   RECT 0.0 331.74 671.84 333.45 ;
   RECT 0.0 333.45 671.84 335.16 ;
   RECT 0.0 335.16 671.84 336.87 ;
   RECT 0.0 336.87 671.84 338.58 ;
   RECT 0.0 338.58 671.84 340.29 ;
   RECT 0.0 340.29 671.84 342.0 ;
   RECT 0.0 342.0 671.84 343.71 ;
   RECT 0.0 343.71 671.84 345.42 ;
   RECT 0.0 345.42 671.84 347.13 ;
   RECT 0.0 347.13 671.84 348.84 ;
   RECT 0.0 348.84 671.84 350.55 ;
   RECT 0.0 350.55 671.84 352.26 ;
   RECT 0.0 352.26 671.84 353.97 ;
   RECT 0.0 353.97 671.84 355.68 ;
   RECT 0.0 355.68 671.84 357.39 ;
   RECT 0.0 357.39 671.84 359.1 ;
   RECT 0.0 359.1 671.84 360.81 ;
   RECT 0.0 360.81 671.84 362.52 ;
   RECT 0.0 362.52 671.84 364.23 ;
   RECT 0.0 364.23 671.84 365.94 ;
   RECT 0.0 365.94 671.84 367.65 ;
   RECT 0.0 367.65 671.84 369.36 ;
   RECT 0.0 369.36 671.84 371.07 ;
   RECT 0.0 371.07 671.84 372.78 ;
   RECT 0.0 372.78 671.84 374.49 ;
   RECT 0.0 374.49 671.84 376.2 ;
   RECT 0.0 376.2 671.84 377.91 ;
   RECT 0.0 377.91 671.84 379.62 ;
   RECT 0.0 379.62 671.84 381.33 ;
   RECT 0.0 381.33 671.84 383.04 ;
   RECT 0.0 383.04 671.84 384.75 ;
   RECT 0.0 384.75 671.84 386.46 ;
   RECT 0.0 386.46 671.84 388.17 ;
   RECT 0.0 388.17 671.84 389.88 ;
   RECT 0.0 389.88 671.84 391.59 ;
   RECT 0.0 391.59 671.84 393.3 ;
   RECT 0.0 393.3 671.84 395.01 ;
   RECT 0.0 395.01 671.84 396.72 ;
   RECT 0.0 396.72 671.84 398.43 ;
   RECT 0.0 398.43 671.84 400.14 ;
   RECT 0.0 400.14 671.84 401.85 ;
   RECT 0.0 401.85 671.84 403.56 ;
   RECT 0.0 403.56 671.84 405.27 ;
   RECT 0.0 405.27 671.84 406.98 ;
   RECT 0.0 406.98 671.84 408.69 ;
   RECT 0.0 408.69 671.84 410.4 ;
 END
END block_1829x2160_148

MACRO block_341x369_84
 CLASS BLOCK ;
 FOREIGN block_341x369_84 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 129.58 BY 70.11 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 20.235 126.445 20.805 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 26.695 126.445 27.265 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 6.935 3.325 7.505 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 7.695 3.325 8.265 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 6.175 3.325 6.745 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 9.215 3.325 9.785 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 10.735 3.325 11.305 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 11.495 3.325 12.065 ;
  END
 END o7
 PIN o8
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 12.255 3.325 12.825 ;
  END
 END o8
 PIN o9
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 13.015 3.325 13.585 ;
  END
 END o9
 PIN o10
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 13.395 4.085 13.965 ;
  END
 END o10
 PIN o11
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 13.775 3.325 14.345 ;
  END
 END o11
 PIN o12
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 15.295 3.325 15.865 ;
  END
 END o12
 PIN o13
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 16.055 3.325 16.625 ;
  END
 END o13
 PIN o14
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 16.815 3.325 17.385 ;
  END
 END o14
 PIN o15
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 12.635 4.085 13.205 ;
  END
 END o15
 PIN o16
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 19.855 3.325 20.425 ;
  END
 END o16
 PIN o17
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 20.615 3.325 21.185 ;
  END
 END o17
 PIN o18
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 21.375 3.325 21.945 ;
  END
 END o18
 PIN o19
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 22.135 3.325 22.705 ;
  END
 END o19
 PIN o20
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 22.895 3.325 23.465 ;
  END
 END o20
 PIN o21
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 18.335 3.325 18.905 ;
  END
 END o21
 PIN o22
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 25.935 3.325 26.505 ;
  END
 END o22
 PIN o23
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 26.695 3.325 27.265 ;
  END
 END o23
 PIN o24
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 27.455 3.325 28.025 ;
  END
 END o24
 PIN o25
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 28.975 3.325 29.545 ;
  END
 END o25
 PIN o26
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 29.735 3.325 30.305 ;
  END
 END o26
 PIN o27
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 25.175 3.325 25.745 ;
  END
 END o27
 PIN o28
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 32.015 3.325 32.585 ;
  END
 END o28
 PIN o29
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 33.535 3.325 34.105 ;
  END
 END o29
 PIN o30
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 34.295 3.325 34.865 ;
  END
 END o30
 PIN o31
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 35.055 3.325 35.625 ;
  END
 END o31
 PIN o32
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 35.815 3.325 36.385 ;
  END
 END o32
 PIN o33
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 31.255 3.325 31.825 ;
  END
 END o33
 PIN o34
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 38.095 126.445 38.665 ;
  END
 END o34
 PIN o35
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 38.855 126.445 39.425 ;
  END
 END o35
 PIN o36
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 39.615 126.445 40.185 ;
  END
 END o36
 PIN o37
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 42.655 126.445 43.225 ;
  END
 END o37
 PIN o38
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 29.735 126.445 30.305 ;
  END
 END o38
 PIN o39
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 21.755 126.445 22.325 ;
  END
 END o39
 PIN o40
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 31.255 126.445 31.825 ;
  END
 END o40
 PIN o41
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 32.015 126.445 32.585 ;
  END
 END o41
 PIN o42
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 33.535 126.445 34.105 ;
  END
 END o42
 PIN o43
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 34.295 126.445 34.865 ;
  END
 END o43
 PIN o44
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 35.055 126.445 35.625 ;
  END
 END o44
 PIN o45
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 30.495 126.445 31.065 ;
  END
 END o45
 PIN o46
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 28.975 126.445 29.545 ;
  END
 END o46
 PIN o47
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 41.135 3.325 41.705 ;
  END
 END o47
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 35.815 126.445 36.385 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 43.035 125.685 43.605 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 32.395 125.685 32.965 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 35.435 125.685 36.005 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 36.955 126.445 37.525 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 36.575 125.685 37.145 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 33.915 125.685 34.485 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 30.115 125.685 30.685 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 40.375 3.325 40.945 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 8.455 3.325 9.025 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 25.935 126.445 26.505 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 25.175 126.445 25.745 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 24.415 126.445 24.985 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 34.675 125.685 35.245 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 30.875 125.685 31.445 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 40.755 126.445 41.325 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 27.455 126.445 28.025 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 38.475 125.685 39.045 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 39.995 125.685 40.565 ;
  END
 END i18
 PIN i19
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 39.235 125.685 39.805 ;
  END
 END i19
 PIN i20
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 124.355 40.375 124.925 40.945 ;
  END
 END i20
 PIN i21
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 8.455 126.445 9.025 ;
  END
 END i21
 PIN i22
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 9.215 126.445 9.785 ;
  END
 END i22
 PIN i23
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 10.735 126.445 11.305 ;
  END
 END i23
 PIN i24
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 11.495 126.445 12.065 ;
  END
 END i24
 PIN i25
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 12.255 126.445 12.825 ;
  END
 END i25
 PIN i26
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 13.015 126.445 13.585 ;
  END
 END i26
 PIN i27
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 8.075 125.685 8.645 ;
  END
 END i27
 PIN i28
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 7.695 126.445 8.265 ;
  END
 END i28
 PIN i29
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 7.315 125.685 7.885 ;
  END
 END i29
 PIN i30
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 6.935 126.445 7.505 ;
  END
 END i30
 PIN i31
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 6.555 125.685 7.125 ;
  END
 END i31
 PIN i32
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 13.775 126.445 14.345 ;
  END
 END i32
 PIN i33
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 15.295 126.445 15.865 ;
  END
 END i33
 PIN i34
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 16.055 126.445 16.625 ;
  END
 END i34
 PIN i35
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 16.815 126.445 17.385 ;
  END
 END i35
 OBS
  LAYER metal1 ;
   RECT 0 0 129.58 70.11 ;
  LAYER via1 ;
   RECT 0 0 129.58 70.11 ;
  LAYER metal2 ;
   RECT 0 0 129.58 70.11 ;
  LAYER via2 ;
   RECT 0 0 129.58 70.11 ;
  LAYER metal3 ;
   RECT 0 0 129.58 70.11 ;
  LAYER via3 ;
   RECT 0 0 129.58 70.11 ;
  LAYER metal4 ;
   RECT 0 0 129.58 70.11 ;
 END
END block_341x369_84

MACRO block_779x1467_106
 CLASS BLOCK ;
 FOREIGN block_779x1467_106 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 296.02 BY 278.73 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 108.395 27.265 108.965 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 92.055 27.265 92.625 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 57.475 27.265 58.045 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 41.135 27.265 41.705 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 24.795 27.265 25.365 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 8.455 27.265 9.025 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 252.795 27.265 253.365 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 169.195 27.265 169.765 ;
  END
 END o7
 PIN o8
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 201.875 27.265 202.445 ;
  END
 END o8
 PIN o9
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 236.455 27.265 237.025 ;
  END
 END o9
 PIN o10
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 185.535 27.265 186.105 ;
  END
 END o10
 PIN o11
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 124.735 27.265 125.305 ;
  END
 END o11
 PIN o12
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 269.135 27.265 269.705 ;
  END
 END o12
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 135.755 4.085 136.325 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 152.855 4.085 153.425 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 141.075 4.085 141.645 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 145.445 4.085 146.015 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 148.295 4.085 148.865 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 4.275 136.135 4.845 136.705 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 4.275 135.375 4.845 135.945 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 134.995 4.085 135.565 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 144.685 4.085 145.255 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 157.795 4.085 158.365 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 4.275 152.475 4.845 153.045 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 149.245 4.085 149.815 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 152.095 4.085 152.665 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 154.185 4.085 154.755 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 156.655 4.085 157.225 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 4.275 158.175 4.845 158.745 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 13.015 134.615 13.585 135.185 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 13.015 147.915 13.585 148.485 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 6.745 27.265 7.315 ;
  END
 END i18
 PIN i19
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 23.085 27.265 23.655 ;
  END
 END i19
 PIN i20
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 238.165 27.265 238.735 ;
  END
 END i20
 PIN i21
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 254.505 27.265 255.075 ;
  END
 END i21
 PIN i22
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 270.845 27.265 271.415 ;
  END
 END i22
 PIN i23
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 39.425 27.265 39.995 ;
  END
 END i23
 PIN i24
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 55.765 27.265 56.335 ;
  END
 END i24
 PIN i25
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 90.345 27.265 90.915 ;
  END
 END i25
 PIN i26
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 106.685 27.265 107.255 ;
  END
 END i26
 PIN i27
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 123.025 27.265 123.595 ;
  END
 END i27
 PIN i28
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 170.905 27.265 171.475 ;
  END
 END i28
 PIN i29
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 187.245 27.265 187.815 ;
  END
 END i29
 PIN i30
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 203.585 27.265 204.155 ;
  END
 END i30
 PIN i31
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.455 41.705 28.025 42.275 ;
  END
 END i31
 PIN i32
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 45.695 27.265 46.265 ;
  END
 END i32
 PIN i33
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 49.875 27.265 50.445 ;
  END
 END i33
 PIN i34
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 33.535 27.265 34.105 ;
  END
 END i34
 PIN i35
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.455 108.965 28.025 109.535 ;
  END
 END i35
 PIN i36
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 112.955 27.265 113.525 ;
  END
 END i36
 PIN i37
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 117.135 27.265 117.705 ;
  END
 END i37
 PIN i38
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 121.125 27.265 121.695 ;
  END
 END i38
 PIN i39
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.455 184.965 28.025 185.535 ;
  END
 END i39
 PIN i40
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 180.975 27.265 181.545 ;
  END
 END i40
 PIN i41
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 176.795 27.265 177.365 ;
  END
 END i41
 PIN i42
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 172.805 27.265 173.375 ;
  END
 END i42
 PIN i43
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.455 252.225 28.025 252.795 ;
  END
 END i43
 PIN i44
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 248.235 27.265 248.805 ;
  END
 END i44
 PIN i45
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 244.055 27.265 244.625 ;
  END
 END i45
 PIN i46
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 260.395 27.265 260.965 ;
  END
 END i46
 PIN i47
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 37.525 27.265 38.095 ;
  END
 END i47
 PIN i48
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 104.785 27.265 105.355 ;
  END
 END i48
 PIN i49
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 189.145 27.265 189.715 ;
  END
 END i49
 PIN i50
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 256.405 27.265 256.975 ;
  END
 END i50
 PIN i51
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 18.335 134.615 18.905 135.185 ;
  END
 END i51
 PIN i52
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 18.335 147.915 18.905 148.485 ;
  END
 END i52
 PIN i53
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.455 7.315 28.025 7.885 ;
  END
 END i53
 PIN i54
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.455 23.655 28.025 24.225 ;
  END
 END i54
 PIN i55
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.455 237.595 28.025 238.165 ;
  END
 END i55
 PIN i56
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.455 253.935 28.025 254.505 ;
  END
 END i56
 PIN i57
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.455 270.275 28.025 270.845 ;
  END
 END i57
 PIN i58
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.455 39.995 28.025 40.565 ;
  END
 END i58
 PIN i59
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.455 56.335 28.025 56.905 ;
  END
 END i59
 PIN i60
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.455 90.915 28.025 91.485 ;
  END
 END i60
 PIN i61
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.455 107.255 28.025 107.825 ;
  END
 END i61
 PIN i62
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.455 123.595 28.025 124.165 ;
  END
 END i62
 PIN i63
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.455 170.335 28.025 170.905 ;
  END
 END i63
 PIN i64
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.455 186.675 28.025 187.245 ;
  END
 END i64
 PIN i65
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.455 203.015 28.025 203.585 ;
  END
 END i65
 PIN i66
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 142.215 4.085 142.785 ;
  END
 END i66
 PIN i67
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 4.275 142.595 4.845 143.165 ;
  END
 END i67
 PIN i68
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.215 7.885 28.785 8.455 ;
  END
 END i68
 PIN i69
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.215 24.225 28.785 24.795 ;
  END
 END i69
 PIN i70
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.215 237.025 28.785 237.595 ;
  END
 END i70
 PIN i71
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.215 253.365 28.785 253.935 ;
  END
 END i71
 PIN i72
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.215 269.705 28.785 270.275 ;
  END
 END i72
 PIN i73
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.215 40.565 28.785 41.135 ;
  END
 END i73
 PIN i74
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.215 56.905 28.785 57.475 ;
  END
 END i74
 PIN i75
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.215 91.485 28.785 92.055 ;
  END
 END i75
 PIN i76
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.215 107.825 28.785 108.395 ;
  END
 END i76
 PIN i77
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.215 124.165 28.785 124.735 ;
  END
 END i77
 PIN i78
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.215 169.765 28.785 170.335 ;
  END
 END i78
 PIN i79
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.215 186.105 28.785 186.675 ;
  END
 END i79
 PIN i80
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.215 202.445 28.785 203.015 ;
  END
 END i80
 PIN i81
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 4.275 134.615 4.845 135.185 ;
  END
 END i81
 PIN i82
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 5.415 134.615 5.985 135.185 ;
  END
 END i82
 PIN i83
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 7.315 134.615 7.885 135.185 ;
  END
 END i83
 PIN i84
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 8.835 134.615 9.405 135.185 ;
  END
 END i84
 PIN i85
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 134.615 10.925 135.185 ;
  END
 END i85
 PIN i86
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 12.255 134.615 12.825 135.185 ;
  END
 END i86
 PIN i87
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 4.275 147.915 4.845 148.485 ;
  END
 END i87
 PIN i88
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 5.415 147.915 5.985 148.485 ;
  END
 END i88
 PIN i89
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 7.315 147.915 7.885 148.485 ;
  END
 END i89
 PIN i90
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 8.835 147.915 9.405 148.485 ;
  END
 END i90
 PIN i91
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 147.915 10.925 148.485 ;
  END
 END i91
 PIN i92
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 12.255 147.915 12.825 148.485 ;
  END
 END i92
 OBS
  LAYER metal1 ;
   RECT 23.18 0.0 296.02 1.71 ;
   RECT 23.18 1.71 296.02 3.42 ;
   RECT 23.18 3.42 296.02 5.13 ;
   RECT 23.18 5.13 296.02 6.84 ;
   RECT 23.18 6.84 296.02 8.55 ;
   RECT 23.18 8.55 296.02 10.26 ;
   RECT 23.18 10.26 296.02 11.97 ;
   RECT 23.18 11.97 296.02 13.68 ;
   RECT 23.18 13.68 296.02 15.39 ;
   RECT 23.18 15.39 296.02 17.1 ;
   RECT 23.18 17.1 296.02 18.81 ;
   RECT 23.18 18.81 296.02 20.52 ;
   RECT 23.18 20.52 296.02 22.23 ;
   RECT 23.18 22.23 296.02 23.94 ;
   RECT 23.18 23.94 296.02 25.65 ;
   RECT 23.18 25.65 296.02 27.36 ;
   RECT 23.18 27.36 296.02 29.07 ;
   RECT 23.18 29.07 296.02 30.78 ;
   RECT 23.18 30.78 296.02 32.49 ;
   RECT 23.18 32.49 296.02 34.2 ;
   RECT 23.18 34.2 296.02 35.91 ;
   RECT 23.18 35.91 296.02 37.62 ;
   RECT 23.18 37.62 296.02 39.33 ;
   RECT 23.18 39.33 296.02 41.04 ;
   RECT 23.18 41.04 296.02 42.75 ;
   RECT 23.18 42.75 296.02 44.46 ;
   RECT 23.18 44.46 296.02 46.17 ;
   RECT 23.18 46.17 296.02 47.88 ;
   RECT 23.18 47.88 296.02 49.59 ;
   RECT 23.18 49.59 296.02 51.3 ;
   RECT 23.18 51.3 296.02 53.01 ;
   RECT 23.18 53.01 296.02 54.72 ;
   RECT 23.18 54.72 296.02 56.43 ;
   RECT 23.18 56.43 296.02 58.14 ;
   RECT 23.18 58.14 296.02 59.85 ;
   RECT 23.18 59.85 296.02 61.56 ;
   RECT 23.18 61.56 296.02 63.27 ;
   RECT 23.18 63.27 296.02 64.98 ;
   RECT 23.18 64.98 296.02 66.69 ;
   RECT 23.18 66.69 296.02 68.4 ;
   RECT 23.18 68.4 296.02 70.11 ;
   RECT 23.18 70.11 296.02 71.82 ;
   RECT 23.18 71.82 296.02 73.53 ;
   RECT 23.18 73.53 296.02 75.24 ;
   RECT 23.18 75.24 296.02 76.95 ;
   RECT 23.18 76.95 296.02 78.66 ;
   RECT 23.18 78.66 296.02 80.37 ;
   RECT 23.18 80.37 296.02 82.08 ;
   RECT 23.18 82.08 296.02 83.79 ;
   RECT 23.18 83.79 296.02 85.5 ;
   RECT 23.18 85.5 296.02 87.21 ;
   RECT 23.18 87.21 296.02 88.92 ;
   RECT 23.18 88.92 296.02 90.63 ;
   RECT 23.18 90.63 296.02 92.34 ;
   RECT 23.18 92.34 296.02 94.05 ;
   RECT 23.18 94.05 296.02 95.76 ;
   RECT 23.18 95.76 296.02 97.47 ;
   RECT 23.18 97.47 296.02 99.18 ;
   RECT 23.18 99.18 296.02 100.89 ;
   RECT 23.18 100.89 296.02 102.6 ;
   RECT 23.18 102.6 296.02 104.31 ;
   RECT 23.18 104.31 296.02 106.02 ;
   RECT 23.18 106.02 296.02 107.73 ;
   RECT 23.18 107.73 296.02 109.44 ;
   RECT 23.18 109.44 296.02 111.15 ;
   RECT 23.18 111.15 296.02 112.86 ;
   RECT 23.18 112.86 296.02 114.57 ;
   RECT 23.18 114.57 296.02 116.28 ;
   RECT 23.18 116.28 296.02 117.99 ;
   RECT 23.18 117.99 296.02 119.7 ;
   RECT 23.18 119.7 296.02 121.41 ;
   RECT 23.18 121.41 296.02 123.12 ;
   RECT 23.18 123.12 296.02 124.83 ;
   RECT 23.18 124.83 296.02 126.54 ;
   RECT 23.18 126.54 296.02 128.25 ;
   RECT 23.18 128.25 296.02 129.96 ;
   RECT 23.18 129.96 296.02 131.67 ;
   RECT 23.18 131.67 296.02 133.38 ;
   RECT 0.0 133.38 296.02 135.09 ;
   RECT 0.0 135.09 296.02 136.8 ;
   RECT 0.0 136.8 296.02 138.51 ;
   RECT 0.0 138.51 296.02 140.22 ;
   RECT 0.0 140.22 296.02 141.93 ;
   RECT 0.0 141.93 296.02 143.64 ;
   RECT 0.0 143.64 296.02 145.35 ;
   RECT 0.0 145.35 296.02 147.06 ;
   RECT 0.0 147.06 296.02 148.77 ;
   RECT 0.0 148.77 296.02 150.48 ;
   RECT 0.0 150.48 296.02 152.19 ;
   RECT 0.0 152.19 296.02 153.9 ;
   RECT 0.0 153.9 296.02 155.61 ;
   RECT 0.0 155.61 296.02 157.32 ;
   RECT 0.0 157.32 296.02 159.03 ;
   RECT 0.0 159.03 296.02 160.74 ;
   RECT 0.0 160.74 296.02 162.45 ;
   RECT 23.18 162.45 296.02 164.16 ;
   RECT 23.18 164.16 296.02 165.87 ;
   RECT 23.18 165.87 296.02 167.58 ;
   RECT 23.18 167.58 296.02 169.29 ;
   RECT 23.18 169.29 296.02 171.0 ;
   RECT 23.18 171.0 296.02 172.71 ;
   RECT 23.18 172.71 296.02 174.42 ;
   RECT 23.18 174.42 296.02 176.13 ;
   RECT 23.18 176.13 296.02 177.84 ;
   RECT 23.18 177.84 296.02 179.55 ;
   RECT 23.18 179.55 296.02 181.26 ;
   RECT 23.18 181.26 296.02 182.97 ;
   RECT 23.18 182.97 296.02 184.68 ;
   RECT 23.18 184.68 296.02 186.39 ;
   RECT 23.18 186.39 296.02 188.1 ;
   RECT 23.18 188.1 296.02 189.81 ;
   RECT 23.18 189.81 296.02 191.52 ;
   RECT 23.18 191.52 296.02 193.23 ;
   RECT 23.18 193.23 296.02 194.94 ;
   RECT 23.18 194.94 296.02 196.65 ;
   RECT 23.18 196.65 296.02 198.36 ;
   RECT 23.18 198.36 296.02 200.07 ;
   RECT 23.18 200.07 296.02 201.78 ;
   RECT 23.18 201.78 296.02 203.49 ;
   RECT 23.18 203.49 296.02 205.2 ;
   RECT 23.18 205.2 296.02 206.91 ;
   RECT 23.18 206.91 296.02 208.62 ;
   RECT 23.18 208.62 296.02 210.33 ;
   RECT 23.18 210.33 296.02 212.04 ;
   RECT 23.18 212.04 296.02 213.75 ;
   RECT 23.18 213.75 296.02 215.46 ;
   RECT 23.18 215.46 296.02 217.17 ;
   RECT 23.18 217.17 296.02 218.88 ;
   RECT 23.18 218.88 296.02 220.59 ;
   RECT 23.18 220.59 296.02 222.3 ;
   RECT 23.18 222.3 296.02 224.01 ;
   RECT 23.18 224.01 296.02 225.72 ;
   RECT 23.18 225.72 296.02 227.43 ;
   RECT 23.18 227.43 296.02 229.14 ;
   RECT 23.18 229.14 296.02 230.85 ;
   RECT 23.18 230.85 296.02 232.56 ;
   RECT 23.18 232.56 296.02 234.27 ;
   RECT 23.18 234.27 296.02 235.98 ;
   RECT 23.18 235.98 296.02 237.69 ;
   RECT 23.18 237.69 296.02 239.4 ;
   RECT 23.18 239.4 296.02 241.11 ;
   RECT 23.18 241.11 296.02 242.82 ;
   RECT 23.18 242.82 296.02 244.53 ;
   RECT 23.18 244.53 296.02 246.24 ;
   RECT 23.18 246.24 296.02 247.95 ;
   RECT 23.18 247.95 296.02 249.66 ;
   RECT 23.18 249.66 296.02 251.37 ;
   RECT 23.18 251.37 296.02 253.08 ;
   RECT 23.18 253.08 296.02 254.79 ;
   RECT 23.18 254.79 296.02 256.5 ;
   RECT 23.18 256.5 296.02 258.21 ;
   RECT 23.18 258.21 296.02 259.92 ;
   RECT 23.18 259.92 296.02 261.63 ;
   RECT 23.18 261.63 296.02 263.34 ;
   RECT 23.18 263.34 296.02 265.05 ;
   RECT 23.18 265.05 296.02 266.76 ;
   RECT 23.18 266.76 296.02 268.47 ;
   RECT 23.18 268.47 296.02 270.18 ;
   RECT 23.18 270.18 296.02 271.89 ;
   RECT 23.18 271.89 296.02 273.6 ;
   RECT 23.18 273.6 296.02 275.31 ;
   RECT 23.18 275.31 296.02 277.02 ;
   RECT 23.18 277.02 296.02 278.73 ;
  LAYER via1 ;
   RECT 23.18 0.0 296.02 1.71 ;
   RECT 23.18 1.71 296.02 3.42 ;
   RECT 23.18 3.42 296.02 5.13 ;
   RECT 23.18 5.13 296.02 6.84 ;
   RECT 23.18 6.84 296.02 8.55 ;
   RECT 23.18 8.55 296.02 10.26 ;
   RECT 23.18 10.26 296.02 11.97 ;
   RECT 23.18 11.97 296.02 13.68 ;
   RECT 23.18 13.68 296.02 15.39 ;
   RECT 23.18 15.39 296.02 17.1 ;
   RECT 23.18 17.1 296.02 18.81 ;
   RECT 23.18 18.81 296.02 20.52 ;
   RECT 23.18 20.52 296.02 22.23 ;
   RECT 23.18 22.23 296.02 23.94 ;
   RECT 23.18 23.94 296.02 25.65 ;
   RECT 23.18 25.65 296.02 27.36 ;
   RECT 23.18 27.36 296.02 29.07 ;
   RECT 23.18 29.07 296.02 30.78 ;
   RECT 23.18 30.78 296.02 32.49 ;
   RECT 23.18 32.49 296.02 34.2 ;
   RECT 23.18 34.2 296.02 35.91 ;
   RECT 23.18 35.91 296.02 37.62 ;
   RECT 23.18 37.62 296.02 39.33 ;
   RECT 23.18 39.33 296.02 41.04 ;
   RECT 23.18 41.04 296.02 42.75 ;
   RECT 23.18 42.75 296.02 44.46 ;
   RECT 23.18 44.46 296.02 46.17 ;
   RECT 23.18 46.17 296.02 47.88 ;
   RECT 23.18 47.88 296.02 49.59 ;
   RECT 23.18 49.59 296.02 51.3 ;
   RECT 23.18 51.3 296.02 53.01 ;
   RECT 23.18 53.01 296.02 54.72 ;
   RECT 23.18 54.72 296.02 56.43 ;
   RECT 23.18 56.43 296.02 58.14 ;
   RECT 23.18 58.14 296.02 59.85 ;
   RECT 23.18 59.85 296.02 61.56 ;
   RECT 23.18 61.56 296.02 63.27 ;
   RECT 23.18 63.27 296.02 64.98 ;
   RECT 23.18 64.98 296.02 66.69 ;
   RECT 23.18 66.69 296.02 68.4 ;
   RECT 23.18 68.4 296.02 70.11 ;
   RECT 23.18 70.11 296.02 71.82 ;
   RECT 23.18 71.82 296.02 73.53 ;
   RECT 23.18 73.53 296.02 75.24 ;
   RECT 23.18 75.24 296.02 76.95 ;
   RECT 23.18 76.95 296.02 78.66 ;
   RECT 23.18 78.66 296.02 80.37 ;
   RECT 23.18 80.37 296.02 82.08 ;
   RECT 23.18 82.08 296.02 83.79 ;
   RECT 23.18 83.79 296.02 85.5 ;
   RECT 23.18 85.5 296.02 87.21 ;
   RECT 23.18 87.21 296.02 88.92 ;
   RECT 23.18 88.92 296.02 90.63 ;
   RECT 23.18 90.63 296.02 92.34 ;
   RECT 23.18 92.34 296.02 94.05 ;
   RECT 23.18 94.05 296.02 95.76 ;
   RECT 23.18 95.76 296.02 97.47 ;
   RECT 23.18 97.47 296.02 99.18 ;
   RECT 23.18 99.18 296.02 100.89 ;
   RECT 23.18 100.89 296.02 102.6 ;
   RECT 23.18 102.6 296.02 104.31 ;
   RECT 23.18 104.31 296.02 106.02 ;
   RECT 23.18 106.02 296.02 107.73 ;
   RECT 23.18 107.73 296.02 109.44 ;
   RECT 23.18 109.44 296.02 111.15 ;
   RECT 23.18 111.15 296.02 112.86 ;
   RECT 23.18 112.86 296.02 114.57 ;
   RECT 23.18 114.57 296.02 116.28 ;
   RECT 23.18 116.28 296.02 117.99 ;
   RECT 23.18 117.99 296.02 119.7 ;
   RECT 23.18 119.7 296.02 121.41 ;
   RECT 23.18 121.41 296.02 123.12 ;
   RECT 23.18 123.12 296.02 124.83 ;
   RECT 23.18 124.83 296.02 126.54 ;
   RECT 23.18 126.54 296.02 128.25 ;
   RECT 23.18 128.25 296.02 129.96 ;
   RECT 23.18 129.96 296.02 131.67 ;
   RECT 23.18 131.67 296.02 133.38 ;
   RECT 0.0 133.38 296.02 135.09 ;
   RECT 0.0 135.09 296.02 136.8 ;
   RECT 0.0 136.8 296.02 138.51 ;
   RECT 0.0 138.51 296.02 140.22 ;
   RECT 0.0 140.22 296.02 141.93 ;
   RECT 0.0 141.93 296.02 143.64 ;
   RECT 0.0 143.64 296.02 145.35 ;
   RECT 0.0 145.35 296.02 147.06 ;
   RECT 0.0 147.06 296.02 148.77 ;
   RECT 0.0 148.77 296.02 150.48 ;
   RECT 0.0 150.48 296.02 152.19 ;
   RECT 0.0 152.19 296.02 153.9 ;
   RECT 0.0 153.9 296.02 155.61 ;
   RECT 0.0 155.61 296.02 157.32 ;
   RECT 0.0 157.32 296.02 159.03 ;
   RECT 0.0 159.03 296.02 160.74 ;
   RECT 0.0 160.74 296.02 162.45 ;
   RECT 23.18 162.45 296.02 164.16 ;
   RECT 23.18 164.16 296.02 165.87 ;
   RECT 23.18 165.87 296.02 167.58 ;
   RECT 23.18 167.58 296.02 169.29 ;
   RECT 23.18 169.29 296.02 171.0 ;
   RECT 23.18 171.0 296.02 172.71 ;
   RECT 23.18 172.71 296.02 174.42 ;
   RECT 23.18 174.42 296.02 176.13 ;
   RECT 23.18 176.13 296.02 177.84 ;
   RECT 23.18 177.84 296.02 179.55 ;
   RECT 23.18 179.55 296.02 181.26 ;
   RECT 23.18 181.26 296.02 182.97 ;
   RECT 23.18 182.97 296.02 184.68 ;
   RECT 23.18 184.68 296.02 186.39 ;
   RECT 23.18 186.39 296.02 188.1 ;
   RECT 23.18 188.1 296.02 189.81 ;
   RECT 23.18 189.81 296.02 191.52 ;
   RECT 23.18 191.52 296.02 193.23 ;
   RECT 23.18 193.23 296.02 194.94 ;
   RECT 23.18 194.94 296.02 196.65 ;
   RECT 23.18 196.65 296.02 198.36 ;
   RECT 23.18 198.36 296.02 200.07 ;
   RECT 23.18 200.07 296.02 201.78 ;
   RECT 23.18 201.78 296.02 203.49 ;
   RECT 23.18 203.49 296.02 205.2 ;
   RECT 23.18 205.2 296.02 206.91 ;
   RECT 23.18 206.91 296.02 208.62 ;
   RECT 23.18 208.62 296.02 210.33 ;
   RECT 23.18 210.33 296.02 212.04 ;
   RECT 23.18 212.04 296.02 213.75 ;
   RECT 23.18 213.75 296.02 215.46 ;
   RECT 23.18 215.46 296.02 217.17 ;
   RECT 23.18 217.17 296.02 218.88 ;
   RECT 23.18 218.88 296.02 220.59 ;
   RECT 23.18 220.59 296.02 222.3 ;
   RECT 23.18 222.3 296.02 224.01 ;
   RECT 23.18 224.01 296.02 225.72 ;
   RECT 23.18 225.72 296.02 227.43 ;
   RECT 23.18 227.43 296.02 229.14 ;
   RECT 23.18 229.14 296.02 230.85 ;
   RECT 23.18 230.85 296.02 232.56 ;
   RECT 23.18 232.56 296.02 234.27 ;
   RECT 23.18 234.27 296.02 235.98 ;
   RECT 23.18 235.98 296.02 237.69 ;
   RECT 23.18 237.69 296.02 239.4 ;
   RECT 23.18 239.4 296.02 241.11 ;
   RECT 23.18 241.11 296.02 242.82 ;
   RECT 23.18 242.82 296.02 244.53 ;
   RECT 23.18 244.53 296.02 246.24 ;
   RECT 23.18 246.24 296.02 247.95 ;
   RECT 23.18 247.95 296.02 249.66 ;
   RECT 23.18 249.66 296.02 251.37 ;
   RECT 23.18 251.37 296.02 253.08 ;
   RECT 23.18 253.08 296.02 254.79 ;
   RECT 23.18 254.79 296.02 256.5 ;
   RECT 23.18 256.5 296.02 258.21 ;
   RECT 23.18 258.21 296.02 259.92 ;
   RECT 23.18 259.92 296.02 261.63 ;
   RECT 23.18 261.63 296.02 263.34 ;
   RECT 23.18 263.34 296.02 265.05 ;
   RECT 23.18 265.05 296.02 266.76 ;
   RECT 23.18 266.76 296.02 268.47 ;
   RECT 23.18 268.47 296.02 270.18 ;
   RECT 23.18 270.18 296.02 271.89 ;
   RECT 23.18 271.89 296.02 273.6 ;
   RECT 23.18 273.6 296.02 275.31 ;
   RECT 23.18 275.31 296.02 277.02 ;
   RECT 23.18 277.02 296.02 278.73 ;
  LAYER metal2 ;
   RECT 23.18 0.0 296.02 1.71 ;
   RECT 23.18 1.71 296.02 3.42 ;
   RECT 23.18 3.42 296.02 5.13 ;
   RECT 23.18 5.13 296.02 6.84 ;
   RECT 23.18 6.84 296.02 8.55 ;
   RECT 23.18 8.55 296.02 10.26 ;
   RECT 23.18 10.26 296.02 11.97 ;
   RECT 23.18 11.97 296.02 13.68 ;
   RECT 23.18 13.68 296.02 15.39 ;
   RECT 23.18 15.39 296.02 17.1 ;
   RECT 23.18 17.1 296.02 18.81 ;
   RECT 23.18 18.81 296.02 20.52 ;
   RECT 23.18 20.52 296.02 22.23 ;
   RECT 23.18 22.23 296.02 23.94 ;
   RECT 23.18 23.94 296.02 25.65 ;
   RECT 23.18 25.65 296.02 27.36 ;
   RECT 23.18 27.36 296.02 29.07 ;
   RECT 23.18 29.07 296.02 30.78 ;
   RECT 23.18 30.78 296.02 32.49 ;
   RECT 23.18 32.49 296.02 34.2 ;
   RECT 23.18 34.2 296.02 35.91 ;
   RECT 23.18 35.91 296.02 37.62 ;
   RECT 23.18 37.62 296.02 39.33 ;
   RECT 23.18 39.33 296.02 41.04 ;
   RECT 23.18 41.04 296.02 42.75 ;
   RECT 23.18 42.75 296.02 44.46 ;
   RECT 23.18 44.46 296.02 46.17 ;
   RECT 23.18 46.17 296.02 47.88 ;
   RECT 23.18 47.88 296.02 49.59 ;
   RECT 23.18 49.59 296.02 51.3 ;
   RECT 23.18 51.3 296.02 53.01 ;
   RECT 23.18 53.01 296.02 54.72 ;
   RECT 23.18 54.72 296.02 56.43 ;
   RECT 23.18 56.43 296.02 58.14 ;
   RECT 23.18 58.14 296.02 59.85 ;
   RECT 23.18 59.85 296.02 61.56 ;
   RECT 23.18 61.56 296.02 63.27 ;
   RECT 23.18 63.27 296.02 64.98 ;
   RECT 23.18 64.98 296.02 66.69 ;
   RECT 23.18 66.69 296.02 68.4 ;
   RECT 23.18 68.4 296.02 70.11 ;
   RECT 23.18 70.11 296.02 71.82 ;
   RECT 23.18 71.82 296.02 73.53 ;
   RECT 23.18 73.53 296.02 75.24 ;
   RECT 23.18 75.24 296.02 76.95 ;
   RECT 23.18 76.95 296.02 78.66 ;
   RECT 23.18 78.66 296.02 80.37 ;
   RECT 23.18 80.37 296.02 82.08 ;
   RECT 23.18 82.08 296.02 83.79 ;
   RECT 23.18 83.79 296.02 85.5 ;
   RECT 23.18 85.5 296.02 87.21 ;
   RECT 23.18 87.21 296.02 88.92 ;
   RECT 23.18 88.92 296.02 90.63 ;
   RECT 23.18 90.63 296.02 92.34 ;
   RECT 23.18 92.34 296.02 94.05 ;
   RECT 23.18 94.05 296.02 95.76 ;
   RECT 23.18 95.76 296.02 97.47 ;
   RECT 23.18 97.47 296.02 99.18 ;
   RECT 23.18 99.18 296.02 100.89 ;
   RECT 23.18 100.89 296.02 102.6 ;
   RECT 23.18 102.6 296.02 104.31 ;
   RECT 23.18 104.31 296.02 106.02 ;
   RECT 23.18 106.02 296.02 107.73 ;
   RECT 23.18 107.73 296.02 109.44 ;
   RECT 23.18 109.44 296.02 111.15 ;
   RECT 23.18 111.15 296.02 112.86 ;
   RECT 23.18 112.86 296.02 114.57 ;
   RECT 23.18 114.57 296.02 116.28 ;
   RECT 23.18 116.28 296.02 117.99 ;
   RECT 23.18 117.99 296.02 119.7 ;
   RECT 23.18 119.7 296.02 121.41 ;
   RECT 23.18 121.41 296.02 123.12 ;
   RECT 23.18 123.12 296.02 124.83 ;
   RECT 23.18 124.83 296.02 126.54 ;
   RECT 23.18 126.54 296.02 128.25 ;
   RECT 23.18 128.25 296.02 129.96 ;
   RECT 23.18 129.96 296.02 131.67 ;
   RECT 23.18 131.67 296.02 133.38 ;
   RECT 0.0 133.38 296.02 135.09 ;
   RECT 0.0 135.09 296.02 136.8 ;
   RECT 0.0 136.8 296.02 138.51 ;
   RECT 0.0 138.51 296.02 140.22 ;
   RECT 0.0 140.22 296.02 141.93 ;
   RECT 0.0 141.93 296.02 143.64 ;
   RECT 0.0 143.64 296.02 145.35 ;
   RECT 0.0 145.35 296.02 147.06 ;
   RECT 0.0 147.06 296.02 148.77 ;
   RECT 0.0 148.77 296.02 150.48 ;
   RECT 0.0 150.48 296.02 152.19 ;
   RECT 0.0 152.19 296.02 153.9 ;
   RECT 0.0 153.9 296.02 155.61 ;
   RECT 0.0 155.61 296.02 157.32 ;
   RECT 0.0 157.32 296.02 159.03 ;
   RECT 0.0 159.03 296.02 160.74 ;
   RECT 0.0 160.74 296.02 162.45 ;
   RECT 23.18 162.45 296.02 164.16 ;
   RECT 23.18 164.16 296.02 165.87 ;
   RECT 23.18 165.87 296.02 167.58 ;
   RECT 23.18 167.58 296.02 169.29 ;
   RECT 23.18 169.29 296.02 171.0 ;
   RECT 23.18 171.0 296.02 172.71 ;
   RECT 23.18 172.71 296.02 174.42 ;
   RECT 23.18 174.42 296.02 176.13 ;
   RECT 23.18 176.13 296.02 177.84 ;
   RECT 23.18 177.84 296.02 179.55 ;
   RECT 23.18 179.55 296.02 181.26 ;
   RECT 23.18 181.26 296.02 182.97 ;
   RECT 23.18 182.97 296.02 184.68 ;
   RECT 23.18 184.68 296.02 186.39 ;
   RECT 23.18 186.39 296.02 188.1 ;
   RECT 23.18 188.1 296.02 189.81 ;
   RECT 23.18 189.81 296.02 191.52 ;
   RECT 23.18 191.52 296.02 193.23 ;
   RECT 23.18 193.23 296.02 194.94 ;
   RECT 23.18 194.94 296.02 196.65 ;
   RECT 23.18 196.65 296.02 198.36 ;
   RECT 23.18 198.36 296.02 200.07 ;
   RECT 23.18 200.07 296.02 201.78 ;
   RECT 23.18 201.78 296.02 203.49 ;
   RECT 23.18 203.49 296.02 205.2 ;
   RECT 23.18 205.2 296.02 206.91 ;
   RECT 23.18 206.91 296.02 208.62 ;
   RECT 23.18 208.62 296.02 210.33 ;
   RECT 23.18 210.33 296.02 212.04 ;
   RECT 23.18 212.04 296.02 213.75 ;
   RECT 23.18 213.75 296.02 215.46 ;
   RECT 23.18 215.46 296.02 217.17 ;
   RECT 23.18 217.17 296.02 218.88 ;
   RECT 23.18 218.88 296.02 220.59 ;
   RECT 23.18 220.59 296.02 222.3 ;
   RECT 23.18 222.3 296.02 224.01 ;
   RECT 23.18 224.01 296.02 225.72 ;
   RECT 23.18 225.72 296.02 227.43 ;
   RECT 23.18 227.43 296.02 229.14 ;
   RECT 23.18 229.14 296.02 230.85 ;
   RECT 23.18 230.85 296.02 232.56 ;
   RECT 23.18 232.56 296.02 234.27 ;
   RECT 23.18 234.27 296.02 235.98 ;
   RECT 23.18 235.98 296.02 237.69 ;
   RECT 23.18 237.69 296.02 239.4 ;
   RECT 23.18 239.4 296.02 241.11 ;
   RECT 23.18 241.11 296.02 242.82 ;
   RECT 23.18 242.82 296.02 244.53 ;
   RECT 23.18 244.53 296.02 246.24 ;
   RECT 23.18 246.24 296.02 247.95 ;
   RECT 23.18 247.95 296.02 249.66 ;
   RECT 23.18 249.66 296.02 251.37 ;
   RECT 23.18 251.37 296.02 253.08 ;
   RECT 23.18 253.08 296.02 254.79 ;
   RECT 23.18 254.79 296.02 256.5 ;
   RECT 23.18 256.5 296.02 258.21 ;
   RECT 23.18 258.21 296.02 259.92 ;
   RECT 23.18 259.92 296.02 261.63 ;
   RECT 23.18 261.63 296.02 263.34 ;
   RECT 23.18 263.34 296.02 265.05 ;
   RECT 23.18 265.05 296.02 266.76 ;
   RECT 23.18 266.76 296.02 268.47 ;
   RECT 23.18 268.47 296.02 270.18 ;
   RECT 23.18 270.18 296.02 271.89 ;
   RECT 23.18 271.89 296.02 273.6 ;
   RECT 23.18 273.6 296.02 275.31 ;
   RECT 23.18 275.31 296.02 277.02 ;
   RECT 23.18 277.02 296.02 278.73 ;
  LAYER via2 ;
   RECT 23.18 0.0 296.02 1.71 ;
   RECT 23.18 1.71 296.02 3.42 ;
   RECT 23.18 3.42 296.02 5.13 ;
   RECT 23.18 5.13 296.02 6.84 ;
   RECT 23.18 6.84 296.02 8.55 ;
   RECT 23.18 8.55 296.02 10.26 ;
   RECT 23.18 10.26 296.02 11.97 ;
   RECT 23.18 11.97 296.02 13.68 ;
   RECT 23.18 13.68 296.02 15.39 ;
   RECT 23.18 15.39 296.02 17.1 ;
   RECT 23.18 17.1 296.02 18.81 ;
   RECT 23.18 18.81 296.02 20.52 ;
   RECT 23.18 20.52 296.02 22.23 ;
   RECT 23.18 22.23 296.02 23.94 ;
   RECT 23.18 23.94 296.02 25.65 ;
   RECT 23.18 25.65 296.02 27.36 ;
   RECT 23.18 27.36 296.02 29.07 ;
   RECT 23.18 29.07 296.02 30.78 ;
   RECT 23.18 30.78 296.02 32.49 ;
   RECT 23.18 32.49 296.02 34.2 ;
   RECT 23.18 34.2 296.02 35.91 ;
   RECT 23.18 35.91 296.02 37.62 ;
   RECT 23.18 37.62 296.02 39.33 ;
   RECT 23.18 39.33 296.02 41.04 ;
   RECT 23.18 41.04 296.02 42.75 ;
   RECT 23.18 42.75 296.02 44.46 ;
   RECT 23.18 44.46 296.02 46.17 ;
   RECT 23.18 46.17 296.02 47.88 ;
   RECT 23.18 47.88 296.02 49.59 ;
   RECT 23.18 49.59 296.02 51.3 ;
   RECT 23.18 51.3 296.02 53.01 ;
   RECT 23.18 53.01 296.02 54.72 ;
   RECT 23.18 54.72 296.02 56.43 ;
   RECT 23.18 56.43 296.02 58.14 ;
   RECT 23.18 58.14 296.02 59.85 ;
   RECT 23.18 59.85 296.02 61.56 ;
   RECT 23.18 61.56 296.02 63.27 ;
   RECT 23.18 63.27 296.02 64.98 ;
   RECT 23.18 64.98 296.02 66.69 ;
   RECT 23.18 66.69 296.02 68.4 ;
   RECT 23.18 68.4 296.02 70.11 ;
   RECT 23.18 70.11 296.02 71.82 ;
   RECT 23.18 71.82 296.02 73.53 ;
   RECT 23.18 73.53 296.02 75.24 ;
   RECT 23.18 75.24 296.02 76.95 ;
   RECT 23.18 76.95 296.02 78.66 ;
   RECT 23.18 78.66 296.02 80.37 ;
   RECT 23.18 80.37 296.02 82.08 ;
   RECT 23.18 82.08 296.02 83.79 ;
   RECT 23.18 83.79 296.02 85.5 ;
   RECT 23.18 85.5 296.02 87.21 ;
   RECT 23.18 87.21 296.02 88.92 ;
   RECT 23.18 88.92 296.02 90.63 ;
   RECT 23.18 90.63 296.02 92.34 ;
   RECT 23.18 92.34 296.02 94.05 ;
   RECT 23.18 94.05 296.02 95.76 ;
   RECT 23.18 95.76 296.02 97.47 ;
   RECT 23.18 97.47 296.02 99.18 ;
   RECT 23.18 99.18 296.02 100.89 ;
   RECT 23.18 100.89 296.02 102.6 ;
   RECT 23.18 102.6 296.02 104.31 ;
   RECT 23.18 104.31 296.02 106.02 ;
   RECT 23.18 106.02 296.02 107.73 ;
   RECT 23.18 107.73 296.02 109.44 ;
   RECT 23.18 109.44 296.02 111.15 ;
   RECT 23.18 111.15 296.02 112.86 ;
   RECT 23.18 112.86 296.02 114.57 ;
   RECT 23.18 114.57 296.02 116.28 ;
   RECT 23.18 116.28 296.02 117.99 ;
   RECT 23.18 117.99 296.02 119.7 ;
   RECT 23.18 119.7 296.02 121.41 ;
   RECT 23.18 121.41 296.02 123.12 ;
   RECT 23.18 123.12 296.02 124.83 ;
   RECT 23.18 124.83 296.02 126.54 ;
   RECT 23.18 126.54 296.02 128.25 ;
   RECT 23.18 128.25 296.02 129.96 ;
   RECT 23.18 129.96 296.02 131.67 ;
   RECT 23.18 131.67 296.02 133.38 ;
   RECT 0.0 133.38 296.02 135.09 ;
   RECT 0.0 135.09 296.02 136.8 ;
   RECT 0.0 136.8 296.02 138.51 ;
   RECT 0.0 138.51 296.02 140.22 ;
   RECT 0.0 140.22 296.02 141.93 ;
   RECT 0.0 141.93 296.02 143.64 ;
   RECT 0.0 143.64 296.02 145.35 ;
   RECT 0.0 145.35 296.02 147.06 ;
   RECT 0.0 147.06 296.02 148.77 ;
   RECT 0.0 148.77 296.02 150.48 ;
   RECT 0.0 150.48 296.02 152.19 ;
   RECT 0.0 152.19 296.02 153.9 ;
   RECT 0.0 153.9 296.02 155.61 ;
   RECT 0.0 155.61 296.02 157.32 ;
   RECT 0.0 157.32 296.02 159.03 ;
   RECT 0.0 159.03 296.02 160.74 ;
   RECT 0.0 160.74 296.02 162.45 ;
   RECT 23.18 162.45 296.02 164.16 ;
   RECT 23.18 164.16 296.02 165.87 ;
   RECT 23.18 165.87 296.02 167.58 ;
   RECT 23.18 167.58 296.02 169.29 ;
   RECT 23.18 169.29 296.02 171.0 ;
   RECT 23.18 171.0 296.02 172.71 ;
   RECT 23.18 172.71 296.02 174.42 ;
   RECT 23.18 174.42 296.02 176.13 ;
   RECT 23.18 176.13 296.02 177.84 ;
   RECT 23.18 177.84 296.02 179.55 ;
   RECT 23.18 179.55 296.02 181.26 ;
   RECT 23.18 181.26 296.02 182.97 ;
   RECT 23.18 182.97 296.02 184.68 ;
   RECT 23.18 184.68 296.02 186.39 ;
   RECT 23.18 186.39 296.02 188.1 ;
   RECT 23.18 188.1 296.02 189.81 ;
   RECT 23.18 189.81 296.02 191.52 ;
   RECT 23.18 191.52 296.02 193.23 ;
   RECT 23.18 193.23 296.02 194.94 ;
   RECT 23.18 194.94 296.02 196.65 ;
   RECT 23.18 196.65 296.02 198.36 ;
   RECT 23.18 198.36 296.02 200.07 ;
   RECT 23.18 200.07 296.02 201.78 ;
   RECT 23.18 201.78 296.02 203.49 ;
   RECT 23.18 203.49 296.02 205.2 ;
   RECT 23.18 205.2 296.02 206.91 ;
   RECT 23.18 206.91 296.02 208.62 ;
   RECT 23.18 208.62 296.02 210.33 ;
   RECT 23.18 210.33 296.02 212.04 ;
   RECT 23.18 212.04 296.02 213.75 ;
   RECT 23.18 213.75 296.02 215.46 ;
   RECT 23.18 215.46 296.02 217.17 ;
   RECT 23.18 217.17 296.02 218.88 ;
   RECT 23.18 218.88 296.02 220.59 ;
   RECT 23.18 220.59 296.02 222.3 ;
   RECT 23.18 222.3 296.02 224.01 ;
   RECT 23.18 224.01 296.02 225.72 ;
   RECT 23.18 225.72 296.02 227.43 ;
   RECT 23.18 227.43 296.02 229.14 ;
   RECT 23.18 229.14 296.02 230.85 ;
   RECT 23.18 230.85 296.02 232.56 ;
   RECT 23.18 232.56 296.02 234.27 ;
   RECT 23.18 234.27 296.02 235.98 ;
   RECT 23.18 235.98 296.02 237.69 ;
   RECT 23.18 237.69 296.02 239.4 ;
   RECT 23.18 239.4 296.02 241.11 ;
   RECT 23.18 241.11 296.02 242.82 ;
   RECT 23.18 242.82 296.02 244.53 ;
   RECT 23.18 244.53 296.02 246.24 ;
   RECT 23.18 246.24 296.02 247.95 ;
   RECT 23.18 247.95 296.02 249.66 ;
   RECT 23.18 249.66 296.02 251.37 ;
   RECT 23.18 251.37 296.02 253.08 ;
   RECT 23.18 253.08 296.02 254.79 ;
   RECT 23.18 254.79 296.02 256.5 ;
   RECT 23.18 256.5 296.02 258.21 ;
   RECT 23.18 258.21 296.02 259.92 ;
   RECT 23.18 259.92 296.02 261.63 ;
   RECT 23.18 261.63 296.02 263.34 ;
   RECT 23.18 263.34 296.02 265.05 ;
   RECT 23.18 265.05 296.02 266.76 ;
   RECT 23.18 266.76 296.02 268.47 ;
   RECT 23.18 268.47 296.02 270.18 ;
   RECT 23.18 270.18 296.02 271.89 ;
   RECT 23.18 271.89 296.02 273.6 ;
   RECT 23.18 273.6 296.02 275.31 ;
   RECT 23.18 275.31 296.02 277.02 ;
   RECT 23.18 277.02 296.02 278.73 ;
  LAYER metal3 ;
   RECT 23.18 0.0 296.02 1.71 ;
   RECT 23.18 1.71 296.02 3.42 ;
   RECT 23.18 3.42 296.02 5.13 ;
   RECT 23.18 5.13 296.02 6.84 ;
   RECT 23.18 6.84 296.02 8.55 ;
   RECT 23.18 8.55 296.02 10.26 ;
   RECT 23.18 10.26 296.02 11.97 ;
   RECT 23.18 11.97 296.02 13.68 ;
   RECT 23.18 13.68 296.02 15.39 ;
   RECT 23.18 15.39 296.02 17.1 ;
   RECT 23.18 17.1 296.02 18.81 ;
   RECT 23.18 18.81 296.02 20.52 ;
   RECT 23.18 20.52 296.02 22.23 ;
   RECT 23.18 22.23 296.02 23.94 ;
   RECT 23.18 23.94 296.02 25.65 ;
   RECT 23.18 25.65 296.02 27.36 ;
   RECT 23.18 27.36 296.02 29.07 ;
   RECT 23.18 29.07 296.02 30.78 ;
   RECT 23.18 30.78 296.02 32.49 ;
   RECT 23.18 32.49 296.02 34.2 ;
   RECT 23.18 34.2 296.02 35.91 ;
   RECT 23.18 35.91 296.02 37.62 ;
   RECT 23.18 37.62 296.02 39.33 ;
   RECT 23.18 39.33 296.02 41.04 ;
   RECT 23.18 41.04 296.02 42.75 ;
   RECT 23.18 42.75 296.02 44.46 ;
   RECT 23.18 44.46 296.02 46.17 ;
   RECT 23.18 46.17 296.02 47.88 ;
   RECT 23.18 47.88 296.02 49.59 ;
   RECT 23.18 49.59 296.02 51.3 ;
   RECT 23.18 51.3 296.02 53.01 ;
   RECT 23.18 53.01 296.02 54.72 ;
   RECT 23.18 54.72 296.02 56.43 ;
   RECT 23.18 56.43 296.02 58.14 ;
   RECT 23.18 58.14 296.02 59.85 ;
   RECT 23.18 59.85 296.02 61.56 ;
   RECT 23.18 61.56 296.02 63.27 ;
   RECT 23.18 63.27 296.02 64.98 ;
   RECT 23.18 64.98 296.02 66.69 ;
   RECT 23.18 66.69 296.02 68.4 ;
   RECT 23.18 68.4 296.02 70.11 ;
   RECT 23.18 70.11 296.02 71.82 ;
   RECT 23.18 71.82 296.02 73.53 ;
   RECT 23.18 73.53 296.02 75.24 ;
   RECT 23.18 75.24 296.02 76.95 ;
   RECT 23.18 76.95 296.02 78.66 ;
   RECT 23.18 78.66 296.02 80.37 ;
   RECT 23.18 80.37 296.02 82.08 ;
   RECT 23.18 82.08 296.02 83.79 ;
   RECT 23.18 83.79 296.02 85.5 ;
   RECT 23.18 85.5 296.02 87.21 ;
   RECT 23.18 87.21 296.02 88.92 ;
   RECT 23.18 88.92 296.02 90.63 ;
   RECT 23.18 90.63 296.02 92.34 ;
   RECT 23.18 92.34 296.02 94.05 ;
   RECT 23.18 94.05 296.02 95.76 ;
   RECT 23.18 95.76 296.02 97.47 ;
   RECT 23.18 97.47 296.02 99.18 ;
   RECT 23.18 99.18 296.02 100.89 ;
   RECT 23.18 100.89 296.02 102.6 ;
   RECT 23.18 102.6 296.02 104.31 ;
   RECT 23.18 104.31 296.02 106.02 ;
   RECT 23.18 106.02 296.02 107.73 ;
   RECT 23.18 107.73 296.02 109.44 ;
   RECT 23.18 109.44 296.02 111.15 ;
   RECT 23.18 111.15 296.02 112.86 ;
   RECT 23.18 112.86 296.02 114.57 ;
   RECT 23.18 114.57 296.02 116.28 ;
   RECT 23.18 116.28 296.02 117.99 ;
   RECT 23.18 117.99 296.02 119.7 ;
   RECT 23.18 119.7 296.02 121.41 ;
   RECT 23.18 121.41 296.02 123.12 ;
   RECT 23.18 123.12 296.02 124.83 ;
   RECT 23.18 124.83 296.02 126.54 ;
   RECT 23.18 126.54 296.02 128.25 ;
   RECT 23.18 128.25 296.02 129.96 ;
   RECT 23.18 129.96 296.02 131.67 ;
   RECT 23.18 131.67 296.02 133.38 ;
   RECT 0.0 133.38 296.02 135.09 ;
   RECT 0.0 135.09 296.02 136.8 ;
   RECT 0.0 136.8 296.02 138.51 ;
   RECT 0.0 138.51 296.02 140.22 ;
   RECT 0.0 140.22 296.02 141.93 ;
   RECT 0.0 141.93 296.02 143.64 ;
   RECT 0.0 143.64 296.02 145.35 ;
   RECT 0.0 145.35 296.02 147.06 ;
   RECT 0.0 147.06 296.02 148.77 ;
   RECT 0.0 148.77 296.02 150.48 ;
   RECT 0.0 150.48 296.02 152.19 ;
   RECT 0.0 152.19 296.02 153.9 ;
   RECT 0.0 153.9 296.02 155.61 ;
   RECT 0.0 155.61 296.02 157.32 ;
   RECT 0.0 157.32 296.02 159.03 ;
   RECT 0.0 159.03 296.02 160.74 ;
   RECT 0.0 160.74 296.02 162.45 ;
   RECT 23.18 162.45 296.02 164.16 ;
   RECT 23.18 164.16 296.02 165.87 ;
   RECT 23.18 165.87 296.02 167.58 ;
   RECT 23.18 167.58 296.02 169.29 ;
   RECT 23.18 169.29 296.02 171.0 ;
   RECT 23.18 171.0 296.02 172.71 ;
   RECT 23.18 172.71 296.02 174.42 ;
   RECT 23.18 174.42 296.02 176.13 ;
   RECT 23.18 176.13 296.02 177.84 ;
   RECT 23.18 177.84 296.02 179.55 ;
   RECT 23.18 179.55 296.02 181.26 ;
   RECT 23.18 181.26 296.02 182.97 ;
   RECT 23.18 182.97 296.02 184.68 ;
   RECT 23.18 184.68 296.02 186.39 ;
   RECT 23.18 186.39 296.02 188.1 ;
   RECT 23.18 188.1 296.02 189.81 ;
   RECT 23.18 189.81 296.02 191.52 ;
   RECT 23.18 191.52 296.02 193.23 ;
   RECT 23.18 193.23 296.02 194.94 ;
   RECT 23.18 194.94 296.02 196.65 ;
   RECT 23.18 196.65 296.02 198.36 ;
   RECT 23.18 198.36 296.02 200.07 ;
   RECT 23.18 200.07 296.02 201.78 ;
   RECT 23.18 201.78 296.02 203.49 ;
   RECT 23.18 203.49 296.02 205.2 ;
   RECT 23.18 205.2 296.02 206.91 ;
   RECT 23.18 206.91 296.02 208.62 ;
   RECT 23.18 208.62 296.02 210.33 ;
   RECT 23.18 210.33 296.02 212.04 ;
   RECT 23.18 212.04 296.02 213.75 ;
   RECT 23.18 213.75 296.02 215.46 ;
   RECT 23.18 215.46 296.02 217.17 ;
   RECT 23.18 217.17 296.02 218.88 ;
   RECT 23.18 218.88 296.02 220.59 ;
   RECT 23.18 220.59 296.02 222.3 ;
   RECT 23.18 222.3 296.02 224.01 ;
   RECT 23.18 224.01 296.02 225.72 ;
   RECT 23.18 225.72 296.02 227.43 ;
   RECT 23.18 227.43 296.02 229.14 ;
   RECT 23.18 229.14 296.02 230.85 ;
   RECT 23.18 230.85 296.02 232.56 ;
   RECT 23.18 232.56 296.02 234.27 ;
   RECT 23.18 234.27 296.02 235.98 ;
   RECT 23.18 235.98 296.02 237.69 ;
   RECT 23.18 237.69 296.02 239.4 ;
   RECT 23.18 239.4 296.02 241.11 ;
   RECT 23.18 241.11 296.02 242.82 ;
   RECT 23.18 242.82 296.02 244.53 ;
   RECT 23.18 244.53 296.02 246.24 ;
   RECT 23.18 246.24 296.02 247.95 ;
   RECT 23.18 247.95 296.02 249.66 ;
   RECT 23.18 249.66 296.02 251.37 ;
   RECT 23.18 251.37 296.02 253.08 ;
   RECT 23.18 253.08 296.02 254.79 ;
   RECT 23.18 254.79 296.02 256.5 ;
   RECT 23.18 256.5 296.02 258.21 ;
   RECT 23.18 258.21 296.02 259.92 ;
   RECT 23.18 259.92 296.02 261.63 ;
   RECT 23.18 261.63 296.02 263.34 ;
   RECT 23.18 263.34 296.02 265.05 ;
   RECT 23.18 265.05 296.02 266.76 ;
   RECT 23.18 266.76 296.02 268.47 ;
   RECT 23.18 268.47 296.02 270.18 ;
   RECT 23.18 270.18 296.02 271.89 ;
   RECT 23.18 271.89 296.02 273.6 ;
   RECT 23.18 273.6 296.02 275.31 ;
   RECT 23.18 275.31 296.02 277.02 ;
   RECT 23.18 277.02 296.02 278.73 ;
  LAYER via3 ;
   RECT 23.18 0.0 296.02 1.71 ;
   RECT 23.18 1.71 296.02 3.42 ;
   RECT 23.18 3.42 296.02 5.13 ;
   RECT 23.18 5.13 296.02 6.84 ;
   RECT 23.18 6.84 296.02 8.55 ;
   RECT 23.18 8.55 296.02 10.26 ;
   RECT 23.18 10.26 296.02 11.97 ;
   RECT 23.18 11.97 296.02 13.68 ;
   RECT 23.18 13.68 296.02 15.39 ;
   RECT 23.18 15.39 296.02 17.1 ;
   RECT 23.18 17.1 296.02 18.81 ;
   RECT 23.18 18.81 296.02 20.52 ;
   RECT 23.18 20.52 296.02 22.23 ;
   RECT 23.18 22.23 296.02 23.94 ;
   RECT 23.18 23.94 296.02 25.65 ;
   RECT 23.18 25.65 296.02 27.36 ;
   RECT 23.18 27.36 296.02 29.07 ;
   RECT 23.18 29.07 296.02 30.78 ;
   RECT 23.18 30.78 296.02 32.49 ;
   RECT 23.18 32.49 296.02 34.2 ;
   RECT 23.18 34.2 296.02 35.91 ;
   RECT 23.18 35.91 296.02 37.62 ;
   RECT 23.18 37.62 296.02 39.33 ;
   RECT 23.18 39.33 296.02 41.04 ;
   RECT 23.18 41.04 296.02 42.75 ;
   RECT 23.18 42.75 296.02 44.46 ;
   RECT 23.18 44.46 296.02 46.17 ;
   RECT 23.18 46.17 296.02 47.88 ;
   RECT 23.18 47.88 296.02 49.59 ;
   RECT 23.18 49.59 296.02 51.3 ;
   RECT 23.18 51.3 296.02 53.01 ;
   RECT 23.18 53.01 296.02 54.72 ;
   RECT 23.18 54.72 296.02 56.43 ;
   RECT 23.18 56.43 296.02 58.14 ;
   RECT 23.18 58.14 296.02 59.85 ;
   RECT 23.18 59.85 296.02 61.56 ;
   RECT 23.18 61.56 296.02 63.27 ;
   RECT 23.18 63.27 296.02 64.98 ;
   RECT 23.18 64.98 296.02 66.69 ;
   RECT 23.18 66.69 296.02 68.4 ;
   RECT 23.18 68.4 296.02 70.11 ;
   RECT 23.18 70.11 296.02 71.82 ;
   RECT 23.18 71.82 296.02 73.53 ;
   RECT 23.18 73.53 296.02 75.24 ;
   RECT 23.18 75.24 296.02 76.95 ;
   RECT 23.18 76.95 296.02 78.66 ;
   RECT 23.18 78.66 296.02 80.37 ;
   RECT 23.18 80.37 296.02 82.08 ;
   RECT 23.18 82.08 296.02 83.79 ;
   RECT 23.18 83.79 296.02 85.5 ;
   RECT 23.18 85.5 296.02 87.21 ;
   RECT 23.18 87.21 296.02 88.92 ;
   RECT 23.18 88.92 296.02 90.63 ;
   RECT 23.18 90.63 296.02 92.34 ;
   RECT 23.18 92.34 296.02 94.05 ;
   RECT 23.18 94.05 296.02 95.76 ;
   RECT 23.18 95.76 296.02 97.47 ;
   RECT 23.18 97.47 296.02 99.18 ;
   RECT 23.18 99.18 296.02 100.89 ;
   RECT 23.18 100.89 296.02 102.6 ;
   RECT 23.18 102.6 296.02 104.31 ;
   RECT 23.18 104.31 296.02 106.02 ;
   RECT 23.18 106.02 296.02 107.73 ;
   RECT 23.18 107.73 296.02 109.44 ;
   RECT 23.18 109.44 296.02 111.15 ;
   RECT 23.18 111.15 296.02 112.86 ;
   RECT 23.18 112.86 296.02 114.57 ;
   RECT 23.18 114.57 296.02 116.28 ;
   RECT 23.18 116.28 296.02 117.99 ;
   RECT 23.18 117.99 296.02 119.7 ;
   RECT 23.18 119.7 296.02 121.41 ;
   RECT 23.18 121.41 296.02 123.12 ;
   RECT 23.18 123.12 296.02 124.83 ;
   RECT 23.18 124.83 296.02 126.54 ;
   RECT 23.18 126.54 296.02 128.25 ;
   RECT 23.18 128.25 296.02 129.96 ;
   RECT 23.18 129.96 296.02 131.67 ;
   RECT 23.18 131.67 296.02 133.38 ;
   RECT 0.0 133.38 296.02 135.09 ;
   RECT 0.0 135.09 296.02 136.8 ;
   RECT 0.0 136.8 296.02 138.51 ;
   RECT 0.0 138.51 296.02 140.22 ;
   RECT 0.0 140.22 296.02 141.93 ;
   RECT 0.0 141.93 296.02 143.64 ;
   RECT 0.0 143.64 296.02 145.35 ;
   RECT 0.0 145.35 296.02 147.06 ;
   RECT 0.0 147.06 296.02 148.77 ;
   RECT 0.0 148.77 296.02 150.48 ;
   RECT 0.0 150.48 296.02 152.19 ;
   RECT 0.0 152.19 296.02 153.9 ;
   RECT 0.0 153.9 296.02 155.61 ;
   RECT 0.0 155.61 296.02 157.32 ;
   RECT 0.0 157.32 296.02 159.03 ;
   RECT 0.0 159.03 296.02 160.74 ;
   RECT 0.0 160.74 296.02 162.45 ;
   RECT 23.18 162.45 296.02 164.16 ;
   RECT 23.18 164.16 296.02 165.87 ;
   RECT 23.18 165.87 296.02 167.58 ;
   RECT 23.18 167.58 296.02 169.29 ;
   RECT 23.18 169.29 296.02 171.0 ;
   RECT 23.18 171.0 296.02 172.71 ;
   RECT 23.18 172.71 296.02 174.42 ;
   RECT 23.18 174.42 296.02 176.13 ;
   RECT 23.18 176.13 296.02 177.84 ;
   RECT 23.18 177.84 296.02 179.55 ;
   RECT 23.18 179.55 296.02 181.26 ;
   RECT 23.18 181.26 296.02 182.97 ;
   RECT 23.18 182.97 296.02 184.68 ;
   RECT 23.18 184.68 296.02 186.39 ;
   RECT 23.18 186.39 296.02 188.1 ;
   RECT 23.18 188.1 296.02 189.81 ;
   RECT 23.18 189.81 296.02 191.52 ;
   RECT 23.18 191.52 296.02 193.23 ;
   RECT 23.18 193.23 296.02 194.94 ;
   RECT 23.18 194.94 296.02 196.65 ;
   RECT 23.18 196.65 296.02 198.36 ;
   RECT 23.18 198.36 296.02 200.07 ;
   RECT 23.18 200.07 296.02 201.78 ;
   RECT 23.18 201.78 296.02 203.49 ;
   RECT 23.18 203.49 296.02 205.2 ;
   RECT 23.18 205.2 296.02 206.91 ;
   RECT 23.18 206.91 296.02 208.62 ;
   RECT 23.18 208.62 296.02 210.33 ;
   RECT 23.18 210.33 296.02 212.04 ;
   RECT 23.18 212.04 296.02 213.75 ;
   RECT 23.18 213.75 296.02 215.46 ;
   RECT 23.18 215.46 296.02 217.17 ;
   RECT 23.18 217.17 296.02 218.88 ;
   RECT 23.18 218.88 296.02 220.59 ;
   RECT 23.18 220.59 296.02 222.3 ;
   RECT 23.18 222.3 296.02 224.01 ;
   RECT 23.18 224.01 296.02 225.72 ;
   RECT 23.18 225.72 296.02 227.43 ;
   RECT 23.18 227.43 296.02 229.14 ;
   RECT 23.18 229.14 296.02 230.85 ;
   RECT 23.18 230.85 296.02 232.56 ;
   RECT 23.18 232.56 296.02 234.27 ;
   RECT 23.18 234.27 296.02 235.98 ;
   RECT 23.18 235.98 296.02 237.69 ;
   RECT 23.18 237.69 296.02 239.4 ;
   RECT 23.18 239.4 296.02 241.11 ;
   RECT 23.18 241.11 296.02 242.82 ;
   RECT 23.18 242.82 296.02 244.53 ;
   RECT 23.18 244.53 296.02 246.24 ;
   RECT 23.18 246.24 296.02 247.95 ;
   RECT 23.18 247.95 296.02 249.66 ;
   RECT 23.18 249.66 296.02 251.37 ;
   RECT 23.18 251.37 296.02 253.08 ;
   RECT 23.18 253.08 296.02 254.79 ;
   RECT 23.18 254.79 296.02 256.5 ;
   RECT 23.18 256.5 296.02 258.21 ;
   RECT 23.18 258.21 296.02 259.92 ;
   RECT 23.18 259.92 296.02 261.63 ;
   RECT 23.18 261.63 296.02 263.34 ;
   RECT 23.18 263.34 296.02 265.05 ;
   RECT 23.18 265.05 296.02 266.76 ;
   RECT 23.18 266.76 296.02 268.47 ;
   RECT 23.18 268.47 296.02 270.18 ;
   RECT 23.18 270.18 296.02 271.89 ;
   RECT 23.18 271.89 296.02 273.6 ;
   RECT 23.18 273.6 296.02 275.31 ;
   RECT 23.18 275.31 296.02 277.02 ;
   RECT 23.18 277.02 296.02 278.73 ;
  LAYER metal4 ;
   RECT 23.18 0.0 296.02 1.71 ;
   RECT 23.18 1.71 296.02 3.42 ;
   RECT 23.18 3.42 296.02 5.13 ;
   RECT 23.18 5.13 296.02 6.84 ;
   RECT 23.18 6.84 296.02 8.55 ;
   RECT 23.18 8.55 296.02 10.26 ;
   RECT 23.18 10.26 296.02 11.97 ;
   RECT 23.18 11.97 296.02 13.68 ;
   RECT 23.18 13.68 296.02 15.39 ;
   RECT 23.18 15.39 296.02 17.1 ;
   RECT 23.18 17.1 296.02 18.81 ;
   RECT 23.18 18.81 296.02 20.52 ;
   RECT 23.18 20.52 296.02 22.23 ;
   RECT 23.18 22.23 296.02 23.94 ;
   RECT 23.18 23.94 296.02 25.65 ;
   RECT 23.18 25.65 296.02 27.36 ;
   RECT 23.18 27.36 296.02 29.07 ;
   RECT 23.18 29.07 296.02 30.78 ;
   RECT 23.18 30.78 296.02 32.49 ;
   RECT 23.18 32.49 296.02 34.2 ;
   RECT 23.18 34.2 296.02 35.91 ;
   RECT 23.18 35.91 296.02 37.62 ;
   RECT 23.18 37.62 296.02 39.33 ;
   RECT 23.18 39.33 296.02 41.04 ;
   RECT 23.18 41.04 296.02 42.75 ;
   RECT 23.18 42.75 296.02 44.46 ;
   RECT 23.18 44.46 296.02 46.17 ;
   RECT 23.18 46.17 296.02 47.88 ;
   RECT 23.18 47.88 296.02 49.59 ;
   RECT 23.18 49.59 296.02 51.3 ;
   RECT 23.18 51.3 296.02 53.01 ;
   RECT 23.18 53.01 296.02 54.72 ;
   RECT 23.18 54.72 296.02 56.43 ;
   RECT 23.18 56.43 296.02 58.14 ;
   RECT 23.18 58.14 296.02 59.85 ;
   RECT 23.18 59.85 296.02 61.56 ;
   RECT 23.18 61.56 296.02 63.27 ;
   RECT 23.18 63.27 296.02 64.98 ;
   RECT 23.18 64.98 296.02 66.69 ;
   RECT 23.18 66.69 296.02 68.4 ;
   RECT 23.18 68.4 296.02 70.11 ;
   RECT 23.18 70.11 296.02 71.82 ;
   RECT 23.18 71.82 296.02 73.53 ;
   RECT 23.18 73.53 296.02 75.24 ;
   RECT 23.18 75.24 296.02 76.95 ;
   RECT 23.18 76.95 296.02 78.66 ;
   RECT 23.18 78.66 296.02 80.37 ;
   RECT 23.18 80.37 296.02 82.08 ;
   RECT 23.18 82.08 296.02 83.79 ;
   RECT 23.18 83.79 296.02 85.5 ;
   RECT 23.18 85.5 296.02 87.21 ;
   RECT 23.18 87.21 296.02 88.92 ;
   RECT 23.18 88.92 296.02 90.63 ;
   RECT 23.18 90.63 296.02 92.34 ;
   RECT 23.18 92.34 296.02 94.05 ;
   RECT 23.18 94.05 296.02 95.76 ;
   RECT 23.18 95.76 296.02 97.47 ;
   RECT 23.18 97.47 296.02 99.18 ;
   RECT 23.18 99.18 296.02 100.89 ;
   RECT 23.18 100.89 296.02 102.6 ;
   RECT 23.18 102.6 296.02 104.31 ;
   RECT 23.18 104.31 296.02 106.02 ;
   RECT 23.18 106.02 296.02 107.73 ;
   RECT 23.18 107.73 296.02 109.44 ;
   RECT 23.18 109.44 296.02 111.15 ;
   RECT 23.18 111.15 296.02 112.86 ;
   RECT 23.18 112.86 296.02 114.57 ;
   RECT 23.18 114.57 296.02 116.28 ;
   RECT 23.18 116.28 296.02 117.99 ;
   RECT 23.18 117.99 296.02 119.7 ;
   RECT 23.18 119.7 296.02 121.41 ;
   RECT 23.18 121.41 296.02 123.12 ;
   RECT 23.18 123.12 296.02 124.83 ;
   RECT 23.18 124.83 296.02 126.54 ;
   RECT 23.18 126.54 296.02 128.25 ;
   RECT 23.18 128.25 296.02 129.96 ;
   RECT 23.18 129.96 296.02 131.67 ;
   RECT 23.18 131.67 296.02 133.38 ;
   RECT 0.0 133.38 296.02 135.09 ;
   RECT 0.0 135.09 296.02 136.8 ;
   RECT 0.0 136.8 296.02 138.51 ;
   RECT 0.0 138.51 296.02 140.22 ;
   RECT 0.0 140.22 296.02 141.93 ;
   RECT 0.0 141.93 296.02 143.64 ;
   RECT 0.0 143.64 296.02 145.35 ;
   RECT 0.0 145.35 296.02 147.06 ;
   RECT 0.0 147.06 296.02 148.77 ;
   RECT 0.0 148.77 296.02 150.48 ;
   RECT 0.0 150.48 296.02 152.19 ;
   RECT 0.0 152.19 296.02 153.9 ;
   RECT 0.0 153.9 296.02 155.61 ;
   RECT 0.0 155.61 296.02 157.32 ;
   RECT 0.0 157.32 296.02 159.03 ;
   RECT 0.0 159.03 296.02 160.74 ;
   RECT 0.0 160.74 296.02 162.45 ;
   RECT 23.18 162.45 296.02 164.16 ;
   RECT 23.18 164.16 296.02 165.87 ;
   RECT 23.18 165.87 296.02 167.58 ;
   RECT 23.18 167.58 296.02 169.29 ;
   RECT 23.18 169.29 296.02 171.0 ;
   RECT 23.18 171.0 296.02 172.71 ;
   RECT 23.18 172.71 296.02 174.42 ;
   RECT 23.18 174.42 296.02 176.13 ;
   RECT 23.18 176.13 296.02 177.84 ;
   RECT 23.18 177.84 296.02 179.55 ;
   RECT 23.18 179.55 296.02 181.26 ;
   RECT 23.18 181.26 296.02 182.97 ;
   RECT 23.18 182.97 296.02 184.68 ;
   RECT 23.18 184.68 296.02 186.39 ;
   RECT 23.18 186.39 296.02 188.1 ;
   RECT 23.18 188.1 296.02 189.81 ;
   RECT 23.18 189.81 296.02 191.52 ;
   RECT 23.18 191.52 296.02 193.23 ;
   RECT 23.18 193.23 296.02 194.94 ;
   RECT 23.18 194.94 296.02 196.65 ;
   RECT 23.18 196.65 296.02 198.36 ;
   RECT 23.18 198.36 296.02 200.07 ;
   RECT 23.18 200.07 296.02 201.78 ;
   RECT 23.18 201.78 296.02 203.49 ;
   RECT 23.18 203.49 296.02 205.2 ;
   RECT 23.18 205.2 296.02 206.91 ;
   RECT 23.18 206.91 296.02 208.62 ;
   RECT 23.18 208.62 296.02 210.33 ;
   RECT 23.18 210.33 296.02 212.04 ;
   RECT 23.18 212.04 296.02 213.75 ;
   RECT 23.18 213.75 296.02 215.46 ;
   RECT 23.18 215.46 296.02 217.17 ;
   RECT 23.18 217.17 296.02 218.88 ;
   RECT 23.18 218.88 296.02 220.59 ;
   RECT 23.18 220.59 296.02 222.3 ;
   RECT 23.18 222.3 296.02 224.01 ;
   RECT 23.18 224.01 296.02 225.72 ;
   RECT 23.18 225.72 296.02 227.43 ;
   RECT 23.18 227.43 296.02 229.14 ;
   RECT 23.18 229.14 296.02 230.85 ;
   RECT 23.18 230.85 296.02 232.56 ;
   RECT 23.18 232.56 296.02 234.27 ;
   RECT 23.18 234.27 296.02 235.98 ;
   RECT 23.18 235.98 296.02 237.69 ;
   RECT 23.18 237.69 296.02 239.4 ;
   RECT 23.18 239.4 296.02 241.11 ;
   RECT 23.18 241.11 296.02 242.82 ;
   RECT 23.18 242.82 296.02 244.53 ;
   RECT 23.18 244.53 296.02 246.24 ;
   RECT 23.18 246.24 296.02 247.95 ;
   RECT 23.18 247.95 296.02 249.66 ;
   RECT 23.18 249.66 296.02 251.37 ;
   RECT 23.18 251.37 296.02 253.08 ;
   RECT 23.18 253.08 296.02 254.79 ;
   RECT 23.18 254.79 296.02 256.5 ;
   RECT 23.18 256.5 296.02 258.21 ;
   RECT 23.18 258.21 296.02 259.92 ;
   RECT 23.18 259.92 296.02 261.63 ;
   RECT 23.18 261.63 296.02 263.34 ;
   RECT 23.18 263.34 296.02 265.05 ;
   RECT 23.18 265.05 296.02 266.76 ;
   RECT 23.18 266.76 296.02 268.47 ;
   RECT 23.18 268.47 296.02 270.18 ;
   RECT 23.18 270.18 296.02 271.89 ;
   RECT 23.18 271.89 296.02 273.6 ;
   RECT 23.18 273.6 296.02 275.31 ;
   RECT 23.18 275.31 296.02 277.02 ;
   RECT 23.18 277.02 296.02 278.73 ;
 END
END block_779x1467_106

MACRO block_1829x2502_263
 CLASS BLOCK ;
 FOREIGN block_1829x2502_263 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 695.02 BY 475.38 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 469.585 26.885 470.155 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 461.415 26.885 461.985 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 387.885 26.885 388.455 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 379.715 26.885 380.285 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 371.545 26.885 372.115 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 345.135 26.885 345.705 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 336.965 26.885 337.535 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 328.795 26.885 329.365 ;
  END
 END o7
 PIN o8
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 320.625 26.885 321.195 ;
  END
 END o8
 PIN o9
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 312.455 26.885 313.025 ;
  END
 END o9
 PIN o10
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 304.285 26.885 304.855 ;
  END
 END o10
 PIN o11
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 296.115 26.885 296.685 ;
  END
 END o11
 PIN o12
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 453.245 26.885 453.815 ;
  END
 END o12
 PIN o13
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 287.945 26.885 288.515 ;
  END
 END o13
 PIN o14
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 279.775 26.885 280.345 ;
  END
 END o14
 PIN o15
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 271.605 26.885 272.175 ;
  END
 END o15
 PIN o16
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 263.435 26.885 264.005 ;
  END
 END o16
 PIN o17
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 255.265 26.885 255.835 ;
  END
 END o17
 PIN o18
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 247.095 26.885 247.665 ;
  END
 END o18
 PIN o19
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 210.615 26.885 211.185 ;
  END
 END o19
 PIN o20
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 202.445 26.885 203.015 ;
  END
 END o20
 PIN o21
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 194.275 26.885 194.845 ;
  END
 END o21
 PIN o22
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 186.105 26.885 186.675 ;
  END
 END o22
 PIN o23
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 445.075 26.885 445.645 ;
  END
 END o23
 PIN o24
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 177.935 26.885 178.505 ;
  END
 END o24
 PIN o25
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 169.765 26.885 170.335 ;
  END
 END o25
 PIN o26
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 161.595 26.885 162.165 ;
  END
 END o26
 PIN o27
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 153.425 26.885 153.995 ;
  END
 END o27
 PIN o28
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 145.255 26.885 145.825 ;
  END
 END o28
 PIN o29
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 137.085 26.885 137.655 ;
  END
 END o29
 PIN o30
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 128.915 26.885 129.485 ;
  END
 END o30
 PIN o31
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 120.745 26.885 121.315 ;
  END
 END o31
 PIN o32
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 94.335 26.885 94.905 ;
  END
 END o32
 PIN o33
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 86.165 26.885 86.735 ;
  END
 END o33
 PIN o34
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 436.905 26.885 437.475 ;
  END
 END o34
 PIN o35
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 77.995 26.885 78.565 ;
  END
 END o35
 PIN o36
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 69.825 26.885 70.395 ;
  END
 END o36
 PIN o37
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 61.655 26.885 62.225 ;
  END
 END o37
 PIN o38
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 53.485 26.885 54.055 ;
  END
 END o38
 PIN o39
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 45.315 26.885 45.885 ;
  END
 END o39
 PIN o40
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 37.145 26.885 37.715 ;
  END
 END o40
 PIN o41
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 28.975 26.885 29.545 ;
  END
 END o41
 PIN o42
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 20.805 26.885 21.375 ;
  END
 END o42
 PIN o43
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 12.635 26.885 13.205 ;
  END
 END o43
 PIN o44
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 4.465 26.885 5.035 ;
  END
 END o44
 PIN o45
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 428.735 26.885 429.305 ;
  END
 END o45
 PIN o46
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 420.565 26.885 421.135 ;
  END
 END o46
 PIN o47
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 412.395 26.885 412.965 ;
  END
 END o47
 PIN o48
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 404.225 26.885 404.795 ;
  END
 END o48
 PIN o49
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 396.055 26.885 396.625 ;
  END
 END o49
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 240.065 3.705 240.635 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 218.405 3.705 218.975 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 222.965 3.705 223.535 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 234.745 3.705 235.315 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 230.375 3.705 230.945 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 239.685 4.465 240.255 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 240.445 4.465 241.015 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 240.825 3.705 241.395 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 231.135 3.705 231.705 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 218.025 4.465 218.595 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 223.345 4.465 223.915 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 226.575 3.705 227.145 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 219.165 3.705 219.735 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 223.725 3.705 224.295 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 221.635 3.705 222.205 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 218.785 4.465 219.355 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 217.645 3.705 218.215 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 14.155 241.205 14.725 241.775 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 16.055 241.205 16.625 241.775 ;
  END
 END i18
 PIN i19
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 14.155 227.905 14.725 228.475 ;
  END
 END i19
 PIN i20
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 16.055 227.905 16.625 228.475 ;
  END
 END i20
 PIN i21
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 471.295 26.885 471.865 ;
  END
 END i21
 PIN i22
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 463.125 26.885 463.695 ;
  END
 END i22
 PIN i23
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 389.595 26.885 390.165 ;
  END
 END i23
 PIN i24
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 381.425 26.885 381.995 ;
  END
 END i24
 PIN i25
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 373.255 26.885 373.825 ;
  END
 END i25
 PIN i26
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 346.845 26.885 347.415 ;
  END
 END i26
 PIN i27
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 338.675 26.885 339.245 ;
  END
 END i27
 PIN i28
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 330.505 26.885 331.075 ;
  END
 END i28
 PIN i29
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 322.335 26.885 322.905 ;
  END
 END i29
 PIN i30
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 314.165 26.885 314.735 ;
  END
 END i30
 PIN i31
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 305.995 26.885 306.565 ;
  END
 END i31
 PIN i32
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 297.825 26.885 298.395 ;
  END
 END i32
 PIN i33
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 454.955 26.885 455.525 ;
  END
 END i33
 PIN i34
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 289.655 26.885 290.225 ;
  END
 END i34
 PIN i35
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 281.485 26.885 282.055 ;
  END
 END i35
 PIN i36
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 273.315 26.885 273.885 ;
  END
 END i36
 PIN i37
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 265.145 26.885 265.715 ;
  END
 END i37
 PIN i38
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 256.975 26.885 257.545 ;
  END
 END i38
 PIN i39
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 248.805 26.885 249.375 ;
  END
 END i39
 PIN i40
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 208.905 26.885 209.475 ;
  END
 END i40
 PIN i41
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 200.735 26.885 201.305 ;
  END
 END i41
 PIN i42
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 192.565 26.885 193.135 ;
  END
 END i42
 PIN i43
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 184.395 26.885 184.965 ;
  END
 END i43
 PIN i44
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 446.785 26.885 447.355 ;
  END
 END i44
 PIN i45
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 176.225 26.885 176.795 ;
  END
 END i45
 PIN i46
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 168.055 26.885 168.625 ;
  END
 END i46
 PIN i47
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 159.885 26.885 160.455 ;
  END
 END i47
 PIN i48
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 151.715 26.885 152.285 ;
  END
 END i48
 PIN i49
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 143.545 26.885 144.115 ;
  END
 END i49
 PIN i50
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 135.375 26.885 135.945 ;
  END
 END i50
 PIN i51
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 127.205 26.885 127.775 ;
  END
 END i51
 PIN i52
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 119.035 26.885 119.605 ;
  END
 END i52
 PIN i53
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 92.625 26.885 93.195 ;
  END
 END i53
 PIN i54
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 84.455 26.885 85.025 ;
  END
 END i54
 PIN i55
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 438.615 26.885 439.185 ;
  END
 END i55
 PIN i56
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 76.285 26.885 76.855 ;
  END
 END i56
 PIN i57
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 68.115 26.885 68.685 ;
  END
 END i57
 PIN i58
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 59.945 26.885 60.515 ;
  END
 END i58
 PIN i59
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 51.775 26.885 52.345 ;
  END
 END i59
 PIN i60
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 43.605 26.885 44.175 ;
  END
 END i60
 PIN i61
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 35.435 26.885 36.005 ;
  END
 END i61
 PIN i62
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 27.265 26.885 27.835 ;
  END
 END i62
 PIN i63
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 19.095 26.885 19.665 ;
  END
 END i63
 PIN i64
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 10.925 26.885 11.495 ;
  END
 END i64
 PIN i65
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 2.755 26.885 3.325 ;
  END
 END i65
 PIN i66
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 430.445 26.885 431.015 ;
  END
 END i66
 PIN i67
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 422.275 26.885 422.845 ;
  END
 END i67
 PIN i68
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 414.105 26.885 414.675 ;
  END
 END i68
 PIN i69
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 405.935 26.885 406.505 ;
  END
 END i69
 PIN i70
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 397.765 26.885 398.335 ;
  END
 END i70
 PIN i71
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 391.305 26.885 391.875 ;
  END
 END i71
 PIN i72
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 387.315 27.645 387.885 ;
  END
 END i72
 PIN i73
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 383.135 26.885 383.705 ;
  END
 END i73
 PIN i74
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 403.655 27.645 404.225 ;
  END
 END i74
 PIN i75
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 399.475 26.885 400.045 ;
  END
 END i75
 PIN i76
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 324.045 26.885 324.615 ;
  END
 END i76
 PIN i77
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 320.055 27.645 320.625 ;
  END
 END i77
 PIN i78
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 315.875 26.885 316.445 ;
  END
 END i78
 PIN i79
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 311.885 27.645 312.455 ;
  END
 END i79
 PIN i80
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 307.705 26.885 308.275 ;
  END
 END i80
 PIN i81
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 141.835 26.885 142.405 ;
  END
 END i81
 PIN i82
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 145.825 27.645 146.395 ;
  END
 END i82
 PIN i83
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 150.005 26.885 150.575 ;
  END
 END i83
 PIN i84
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 153.995 27.645 154.565 ;
  END
 END i84
 PIN i85
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 158.175 26.885 158.745 ;
  END
 END i85
 PIN i86
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 74.575 26.885 75.145 ;
  END
 END i86
 PIN i87
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 78.565 27.645 79.135 ;
  END
 END i87
 PIN i88
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 82.745 26.885 83.315 ;
  END
 END i88
 PIN i89
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 62.225 27.645 62.795 ;
  END
 END i89
 PIN i90
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 66.405 26.885 66.975 ;
  END
 END i90
 PIN i91
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 395.485 27.645 396.055 ;
  END
 END i91
 PIN i92
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 328.225 27.645 328.795 ;
  END
 END i92
 PIN i93
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 137.655 27.645 138.225 ;
  END
 END i93
 PIN i94
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 70.395 27.645 70.965 ;
  END
 END i94
 PIN i95
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 17.955 241.205 18.525 241.775 ;
  END
 END i95
 PIN i96
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 17.955 227.905 18.525 228.475 ;
  END
 END i96
 PIN i97
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 470.725 27.645 471.295 ;
  END
 END i97
 PIN i98
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 462.555 27.645 463.125 ;
  END
 END i98
 PIN i99
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 389.025 27.645 389.595 ;
  END
 END i99
 PIN i100
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 380.855 27.645 381.425 ;
  END
 END i100
 PIN i101
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 372.685 27.645 373.255 ;
  END
 END i101
 PIN i102
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 346.275 27.645 346.845 ;
  END
 END i102
 PIN i103
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 338.105 27.645 338.675 ;
  END
 END i103
 PIN i104
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 329.935 27.645 330.505 ;
  END
 END i104
 PIN i105
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 321.765 27.645 322.335 ;
  END
 END i105
 PIN i106
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 313.595 27.645 314.165 ;
  END
 END i106
 PIN i107
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 305.425 27.645 305.995 ;
  END
 END i107
 PIN i108
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 297.255 27.645 297.825 ;
  END
 END i108
 PIN i109
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 454.385 27.645 454.955 ;
  END
 END i109
 PIN i110
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 289.085 27.645 289.655 ;
  END
 END i110
 PIN i111
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 280.915 27.645 281.485 ;
  END
 END i111
 PIN i112
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 272.745 27.645 273.315 ;
  END
 END i112
 PIN i113
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 264.575 27.645 265.145 ;
  END
 END i113
 PIN i114
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 256.405 27.645 256.975 ;
  END
 END i114
 PIN i115
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 248.235 27.645 248.805 ;
  END
 END i115
 PIN i116
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 209.475 27.645 210.045 ;
  END
 END i116
 PIN i117
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 201.305 27.645 201.875 ;
  END
 END i117
 PIN i118
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 193.135 27.645 193.705 ;
  END
 END i118
 PIN i119
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 184.965 27.645 185.535 ;
  END
 END i119
 PIN i120
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 446.215 27.645 446.785 ;
  END
 END i120
 PIN i121
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 176.795 27.645 177.365 ;
  END
 END i121
 PIN i122
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 168.625 27.645 169.195 ;
  END
 END i122
 PIN i123
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 160.455 27.645 161.025 ;
  END
 END i123
 PIN i124
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 152.285 27.645 152.855 ;
  END
 END i124
 PIN i125
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 144.115 27.645 144.685 ;
  END
 END i125
 PIN i126
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 135.945 27.645 136.515 ;
  END
 END i126
 PIN i127
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 127.775 27.645 128.345 ;
  END
 END i127
 PIN i128
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 119.605 27.645 120.175 ;
  END
 END i128
 PIN i129
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 93.195 27.645 93.765 ;
  END
 END i129
 PIN i130
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 85.025 27.645 85.595 ;
  END
 END i130
 PIN i131
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 438.045 27.645 438.615 ;
  END
 END i131
 PIN i132
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 76.855 27.645 77.425 ;
  END
 END i132
 PIN i133
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 68.685 27.645 69.255 ;
  END
 END i133
 PIN i134
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 60.515 27.645 61.085 ;
  END
 END i134
 PIN i135
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 52.345 27.645 52.915 ;
  END
 END i135
 PIN i136
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 44.175 27.645 44.745 ;
  END
 END i136
 PIN i137
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 36.005 27.645 36.575 ;
  END
 END i137
 PIN i138
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 27.835 27.645 28.405 ;
  END
 END i138
 PIN i139
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 19.665 27.645 20.235 ;
  END
 END i139
 PIN i140
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 11.495 27.645 12.065 ;
  END
 END i140
 PIN i141
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 3.325 27.645 3.895 ;
  END
 END i141
 PIN i142
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 429.875 27.645 430.445 ;
  END
 END i142
 PIN i143
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 421.705 27.645 422.275 ;
  END
 END i143
 PIN i144
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 413.535 27.645 414.105 ;
  END
 END i144
 PIN i145
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 405.365 27.645 405.935 ;
  END
 END i145
 PIN i146
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 397.195 27.645 397.765 ;
  END
 END i146
 PIN i147
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 233.605 3.705 234.175 ;
  END
 END i147
 PIN i148
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 233.225 4.465 233.795 ;
  END
 END i148
 PIN i149
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 470.155 28.405 470.725 ;
  END
 END i149
 PIN i150
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 461.985 28.405 462.555 ;
  END
 END i150
 PIN i151
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 388.455 28.405 389.025 ;
  END
 END i151
 PIN i152
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 380.285 28.405 380.855 ;
  END
 END i152
 PIN i153
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 372.115 28.405 372.685 ;
  END
 END i153
 PIN i154
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 345.705 28.405 346.275 ;
  END
 END i154
 PIN i155
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 337.535 28.405 338.105 ;
  END
 END i155
 PIN i156
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 329.365 28.405 329.935 ;
  END
 END i156
 PIN i157
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 321.195 28.405 321.765 ;
  END
 END i157
 PIN i158
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 313.025 28.405 313.595 ;
  END
 END i158
 PIN i159
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 304.855 28.405 305.425 ;
  END
 END i159
 PIN i160
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 296.685 28.405 297.255 ;
  END
 END i160
 PIN i161
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 453.815 28.405 454.385 ;
  END
 END i161
 PIN i162
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 288.515 28.405 289.085 ;
  END
 END i162
 PIN i163
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 280.345 28.405 280.915 ;
  END
 END i163
 PIN i164
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 272.175 28.405 272.745 ;
  END
 END i164
 PIN i165
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 264.005 28.405 264.575 ;
  END
 END i165
 PIN i166
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 255.835 28.405 256.405 ;
  END
 END i166
 PIN i167
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 247.665 28.405 248.235 ;
  END
 END i167
 PIN i168
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 210.045 28.405 210.615 ;
  END
 END i168
 PIN i169
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 201.875 28.405 202.445 ;
  END
 END i169
 PIN i170
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 193.705 28.405 194.275 ;
  END
 END i170
 PIN i171
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 185.535 28.405 186.105 ;
  END
 END i171
 PIN i172
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 445.645 28.405 446.215 ;
  END
 END i172
 PIN i173
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 177.365 28.405 177.935 ;
  END
 END i173
 PIN i174
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 169.195 28.405 169.765 ;
  END
 END i174
 PIN i175
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 161.025 28.405 161.595 ;
  END
 END i175
 PIN i176
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 152.855 28.405 153.425 ;
  END
 END i176
 PIN i177
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 144.685 28.405 145.255 ;
  END
 END i177
 PIN i178
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 136.515 28.405 137.085 ;
  END
 END i178
 PIN i179
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 128.345 28.405 128.915 ;
  END
 END i179
 PIN i180
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 120.175 28.405 120.745 ;
  END
 END i180
 PIN i181
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 93.765 28.405 94.335 ;
  END
 END i181
 PIN i182
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 85.595 28.405 86.165 ;
  END
 END i182
 PIN i183
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 437.475 28.405 438.045 ;
  END
 END i183
 PIN i184
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 77.425 28.405 77.995 ;
  END
 END i184
 PIN i185
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 69.255 28.405 69.825 ;
  END
 END i185
 PIN i186
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 61.085 28.405 61.655 ;
  END
 END i186
 PIN i187
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 52.915 28.405 53.485 ;
  END
 END i187
 PIN i188
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 44.745 28.405 45.315 ;
  END
 END i188
 PIN i189
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 36.575 28.405 37.145 ;
  END
 END i189
 PIN i190
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 28.405 28.405 28.975 ;
  END
 END i190
 PIN i191
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 20.235 28.405 20.805 ;
  END
 END i191
 PIN i192
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 12.065 28.405 12.635 ;
  END
 END i192
 PIN i193
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 3.895 28.405 4.465 ;
  END
 END i193
 PIN i194
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 429.305 28.405 429.875 ;
  END
 END i194
 PIN i195
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 421.135 28.405 421.705 ;
  END
 END i195
 PIN i196
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 412.965 28.405 413.535 ;
  END
 END i196
 PIN i197
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 404.795 28.405 405.365 ;
  END
 END i197
 PIN i198
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 396.625 28.405 397.195 ;
  END
 END i198
 PIN i199
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 4.275 241.205 4.845 241.775 ;
  END
 END i199
 PIN i200
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 5.415 241.205 5.985 241.775 ;
  END
 END i200
 PIN i201
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 6.935 241.205 7.505 241.775 ;
  END
 END i201
 PIN i202
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 8.835 241.205 9.405 241.775 ;
  END
 END i202
 PIN i203
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 241.205 10.925 241.775 ;
  END
 END i203
 PIN i204
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 11.875 241.205 12.445 241.775 ;
  END
 END i204
 PIN i205
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 13.015 241.205 13.585 241.775 ;
  END
 END i205
 PIN i206
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 4.275 227.905 4.845 228.475 ;
  END
 END i206
 PIN i207
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 5.415 227.905 5.985 228.475 ;
  END
 END i207
 PIN i208
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 6.935 227.905 7.505 228.475 ;
  END
 END i208
 PIN i209
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 8.835 227.905 9.405 228.475 ;
  END
 END i209
 PIN i210
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 227.905 10.925 228.475 ;
  END
 END i210
 PIN i211
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 11.875 227.905 12.445 228.475 ;
  END
 END i211
 PIN i212
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 13.015 227.905 13.585 228.475 ;
  END
 END i212
 OBS
  LAYER metal1 ;
   RECT 23.18 0.0 695.02 1.71 ;
   RECT 23.18 1.71 695.02 3.42 ;
   RECT 23.18 3.42 695.02 5.13 ;
   RECT 23.18 5.13 695.02 6.84 ;
   RECT 23.18 6.84 695.02 8.55 ;
   RECT 23.18 8.55 695.02 10.26 ;
   RECT 23.18 10.26 695.02 11.97 ;
   RECT 23.18 11.97 695.02 13.68 ;
   RECT 23.18 13.68 695.02 15.39 ;
   RECT 23.18 15.39 695.02 17.1 ;
   RECT 23.18 17.1 695.02 18.81 ;
   RECT 23.18 18.81 695.02 20.52 ;
   RECT 23.18 20.52 695.02 22.23 ;
   RECT 23.18 22.23 695.02 23.94 ;
   RECT 23.18 23.94 695.02 25.65 ;
   RECT 23.18 25.65 695.02 27.36 ;
   RECT 23.18 27.36 695.02 29.07 ;
   RECT 23.18 29.07 695.02 30.78 ;
   RECT 23.18 30.78 695.02 32.49 ;
   RECT 23.18 32.49 695.02 34.2 ;
   RECT 23.18 34.2 695.02 35.91 ;
   RECT 23.18 35.91 695.02 37.62 ;
   RECT 23.18 37.62 695.02 39.33 ;
   RECT 23.18 39.33 695.02 41.04 ;
   RECT 23.18 41.04 695.02 42.75 ;
   RECT 23.18 42.75 695.02 44.46 ;
   RECT 23.18 44.46 695.02 46.17 ;
   RECT 23.18 46.17 695.02 47.88 ;
   RECT 23.18 47.88 695.02 49.59 ;
   RECT 23.18 49.59 695.02 51.3 ;
   RECT 23.18 51.3 695.02 53.01 ;
   RECT 23.18 53.01 695.02 54.72 ;
   RECT 23.18 54.72 695.02 56.43 ;
   RECT 23.18 56.43 695.02 58.14 ;
   RECT 23.18 58.14 695.02 59.85 ;
   RECT 23.18 59.85 695.02 61.56 ;
   RECT 23.18 61.56 695.02 63.27 ;
   RECT 23.18 63.27 695.02 64.98 ;
   RECT 23.18 64.98 695.02 66.69 ;
   RECT 23.18 66.69 695.02 68.4 ;
   RECT 23.18 68.4 695.02 70.11 ;
   RECT 23.18 70.11 695.02 71.82 ;
   RECT 23.18 71.82 695.02 73.53 ;
   RECT 23.18 73.53 695.02 75.24 ;
   RECT 23.18 75.24 695.02 76.95 ;
   RECT 23.18 76.95 695.02 78.66 ;
   RECT 23.18 78.66 695.02 80.37 ;
   RECT 23.18 80.37 695.02 82.08 ;
   RECT 23.18 82.08 695.02 83.79 ;
   RECT 23.18 83.79 695.02 85.5 ;
   RECT 23.18 85.5 695.02 87.21 ;
   RECT 23.18 87.21 695.02 88.92 ;
   RECT 23.18 88.92 695.02 90.63 ;
   RECT 23.18 90.63 695.02 92.34 ;
   RECT 23.18 92.34 695.02 94.05 ;
   RECT 23.18 94.05 695.02 95.76 ;
   RECT 23.18 95.76 695.02 97.47 ;
   RECT 23.18 97.47 695.02 99.18 ;
   RECT 23.18 99.18 695.02 100.89 ;
   RECT 23.18 100.89 695.02 102.6 ;
   RECT 23.18 102.6 695.02 104.31 ;
   RECT 23.18 104.31 695.02 106.02 ;
   RECT 23.18 106.02 695.02 107.73 ;
   RECT 23.18 107.73 695.02 109.44 ;
   RECT 23.18 109.44 695.02 111.15 ;
   RECT 23.18 111.15 695.02 112.86 ;
   RECT 23.18 112.86 695.02 114.57 ;
   RECT 23.18 114.57 695.02 116.28 ;
   RECT 23.18 116.28 695.02 117.99 ;
   RECT 23.18 117.99 695.02 119.7 ;
   RECT 23.18 119.7 695.02 121.41 ;
   RECT 23.18 121.41 695.02 123.12 ;
   RECT 23.18 123.12 695.02 124.83 ;
   RECT 23.18 124.83 695.02 126.54 ;
   RECT 23.18 126.54 695.02 128.25 ;
   RECT 23.18 128.25 695.02 129.96 ;
   RECT 23.18 129.96 695.02 131.67 ;
   RECT 23.18 131.67 695.02 133.38 ;
   RECT 23.18 133.38 695.02 135.09 ;
   RECT 23.18 135.09 695.02 136.8 ;
   RECT 23.18 136.8 695.02 138.51 ;
   RECT 23.18 138.51 695.02 140.22 ;
   RECT 23.18 140.22 695.02 141.93 ;
   RECT 23.18 141.93 695.02 143.64 ;
   RECT 23.18 143.64 695.02 145.35 ;
   RECT 23.18 145.35 695.02 147.06 ;
   RECT 23.18 147.06 695.02 148.77 ;
   RECT 23.18 148.77 695.02 150.48 ;
   RECT 23.18 150.48 695.02 152.19 ;
   RECT 23.18 152.19 695.02 153.9 ;
   RECT 23.18 153.9 695.02 155.61 ;
   RECT 23.18 155.61 695.02 157.32 ;
   RECT 23.18 157.32 695.02 159.03 ;
   RECT 23.18 159.03 695.02 160.74 ;
   RECT 23.18 160.74 695.02 162.45 ;
   RECT 23.18 162.45 695.02 164.16 ;
   RECT 23.18 164.16 695.02 165.87 ;
   RECT 23.18 165.87 695.02 167.58 ;
   RECT 23.18 167.58 695.02 169.29 ;
   RECT 23.18 169.29 695.02 171.0 ;
   RECT 23.18 171.0 695.02 172.71 ;
   RECT 23.18 172.71 695.02 174.42 ;
   RECT 23.18 174.42 695.02 176.13 ;
   RECT 23.18 176.13 695.02 177.84 ;
   RECT 23.18 177.84 695.02 179.55 ;
   RECT 23.18 179.55 695.02 181.26 ;
   RECT 23.18 181.26 695.02 182.97 ;
   RECT 23.18 182.97 695.02 184.68 ;
   RECT 23.18 184.68 695.02 186.39 ;
   RECT 23.18 186.39 695.02 188.1 ;
   RECT 23.18 188.1 695.02 189.81 ;
   RECT 23.18 189.81 695.02 191.52 ;
   RECT 23.18 191.52 695.02 193.23 ;
   RECT 23.18 193.23 695.02 194.94 ;
   RECT 23.18 194.94 695.02 196.65 ;
   RECT 23.18 196.65 695.02 198.36 ;
   RECT 23.18 198.36 695.02 200.07 ;
   RECT 23.18 200.07 695.02 201.78 ;
   RECT 23.18 201.78 695.02 203.49 ;
   RECT 23.18 203.49 695.02 205.2 ;
   RECT 23.18 205.2 695.02 206.91 ;
   RECT 23.18 206.91 695.02 208.62 ;
   RECT 23.18 208.62 695.02 210.33 ;
   RECT 23.18 210.33 695.02 212.04 ;
   RECT 23.18 212.04 695.02 213.75 ;
   RECT 23.18 213.75 695.02 215.46 ;
   RECT 0.0 215.46 695.02 217.17 ;
   RECT 0.0 217.17 695.02 218.88 ;
   RECT 0.0 218.88 695.02 220.59 ;
   RECT 0.0 220.59 695.02 222.3 ;
   RECT 0.0 222.3 695.02 224.01 ;
   RECT 0.0 224.01 695.02 225.72 ;
   RECT 0.0 225.72 695.02 227.43 ;
   RECT 0.0 227.43 695.02 229.14 ;
   RECT 0.0 229.14 695.02 230.85 ;
   RECT 0.0 230.85 695.02 232.56 ;
   RECT 0.0 232.56 695.02 234.27 ;
   RECT 0.0 234.27 695.02 235.98 ;
   RECT 0.0 235.98 695.02 237.69 ;
   RECT 0.0 237.69 695.02 239.4 ;
   RECT 0.0 239.4 695.02 241.11 ;
   RECT 0.0 241.11 695.02 242.82 ;
   RECT 0.0 242.82 695.02 244.53 ;
   RECT 23.18 244.53 695.02 246.24 ;
   RECT 23.18 246.24 695.02 247.95 ;
   RECT 23.18 247.95 695.02 249.66 ;
   RECT 23.18 249.66 695.02 251.37 ;
   RECT 23.18 251.37 695.02 253.08 ;
   RECT 23.18 253.08 695.02 254.79 ;
   RECT 23.18 254.79 695.02 256.5 ;
   RECT 23.18 256.5 695.02 258.21 ;
   RECT 23.18 258.21 695.02 259.92 ;
   RECT 23.18 259.92 695.02 261.63 ;
   RECT 23.18 261.63 695.02 263.34 ;
   RECT 23.18 263.34 695.02 265.05 ;
   RECT 23.18 265.05 695.02 266.76 ;
   RECT 23.18 266.76 695.02 268.47 ;
   RECT 23.18 268.47 695.02 270.18 ;
   RECT 23.18 270.18 695.02 271.89 ;
   RECT 23.18 271.89 695.02 273.6 ;
   RECT 23.18 273.6 695.02 275.31 ;
   RECT 23.18 275.31 695.02 277.02 ;
   RECT 23.18 277.02 695.02 278.73 ;
   RECT 23.18 278.73 695.02 280.44 ;
   RECT 23.18 280.44 695.02 282.15 ;
   RECT 23.18 282.15 695.02 283.86 ;
   RECT 23.18 283.86 695.02 285.57 ;
   RECT 23.18 285.57 695.02 287.28 ;
   RECT 23.18 287.28 695.02 288.99 ;
   RECT 23.18 288.99 695.02 290.7 ;
   RECT 23.18 290.7 695.02 292.41 ;
   RECT 23.18 292.41 695.02 294.12 ;
   RECT 23.18 294.12 695.02 295.83 ;
   RECT 23.18 295.83 695.02 297.54 ;
   RECT 23.18 297.54 695.02 299.25 ;
   RECT 23.18 299.25 695.02 300.96 ;
   RECT 23.18 300.96 695.02 302.67 ;
   RECT 23.18 302.67 695.02 304.38 ;
   RECT 23.18 304.38 695.02 306.09 ;
   RECT 23.18 306.09 695.02 307.8 ;
   RECT 23.18 307.8 695.02 309.51 ;
   RECT 23.18 309.51 695.02 311.22 ;
   RECT 23.18 311.22 695.02 312.93 ;
   RECT 23.18 312.93 695.02 314.64 ;
   RECT 23.18 314.64 695.02 316.35 ;
   RECT 23.18 316.35 695.02 318.06 ;
   RECT 23.18 318.06 695.02 319.77 ;
   RECT 23.18 319.77 695.02 321.48 ;
   RECT 23.18 321.48 695.02 323.19 ;
   RECT 23.18 323.19 695.02 324.9 ;
   RECT 23.18 324.9 695.02 326.61 ;
   RECT 23.18 326.61 695.02 328.32 ;
   RECT 23.18 328.32 695.02 330.03 ;
   RECT 23.18 330.03 695.02 331.74 ;
   RECT 23.18 331.74 695.02 333.45 ;
   RECT 23.18 333.45 695.02 335.16 ;
   RECT 23.18 335.16 695.02 336.87 ;
   RECT 23.18 336.87 695.02 338.58 ;
   RECT 23.18 338.58 695.02 340.29 ;
   RECT 23.18 340.29 695.02 342.0 ;
   RECT 23.18 342.0 695.02 343.71 ;
   RECT 23.18 343.71 695.02 345.42 ;
   RECT 23.18 345.42 695.02 347.13 ;
   RECT 23.18 347.13 695.02 348.84 ;
   RECT 23.18 348.84 695.02 350.55 ;
   RECT 23.18 350.55 695.02 352.26 ;
   RECT 23.18 352.26 695.02 353.97 ;
   RECT 23.18 353.97 695.02 355.68 ;
   RECT 23.18 355.68 695.02 357.39 ;
   RECT 23.18 357.39 695.02 359.1 ;
   RECT 23.18 359.1 695.02 360.81 ;
   RECT 23.18 360.81 695.02 362.52 ;
   RECT 23.18 362.52 695.02 364.23 ;
   RECT 23.18 364.23 695.02 365.94 ;
   RECT 23.18 365.94 695.02 367.65 ;
   RECT 23.18 367.65 695.02 369.36 ;
   RECT 23.18 369.36 695.02 371.07 ;
   RECT 23.18 371.07 695.02 372.78 ;
   RECT 23.18 372.78 695.02 374.49 ;
   RECT 23.18 374.49 695.02 376.2 ;
   RECT 23.18 376.2 695.02 377.91 ;
   RECT 23.18 377.91 695.02 379.62 ;
   RECT 23.18 379.62 695.02 381.33 ;
   RECT 23.18 381.33 695.02 383.04 ;
   RECT 23.18 383.04 695.02 384.75 ;
   RECT 23.18 384.75 695.02 386.46 ;
   RECT 23.18 386.46 695.02 388.17 ;
   RECT 23.18 388.17 695.02 389.88 ;
   RECT 23.18 389.88 695.02 391.59 ;
   RECT 23.18 391.59 695.02 393.3 ;
   RECT 23.18 393.3 695.02 395.01 ;
   RECT 23.18 395.01 695.02 396.72 ;
   RECT 23.18 396.72 695.02 398.43 ;
   RECT 23.18 398.43 695.02 400.14 ;
   RECT 23.18 400.14 695.02 401.85 ;
   RECT 23.18 401.85 695.02 403.56 ;
   RECT 23.18 403.56 695.02 405.27 ;
   RECT 23.18 405.27 695.02 406.98 ;
   RECT 23.18 406.98 695.02 408.69 ;
   RECT 23.18 408.69 695.02 410.4 ;
   RECT 23.18 410.4 695.02 412.11 ;
   RECT 23.18 412.11 695.02 413.82 ;
   RECT 23.18 413.82 695.02 415.53 ;
   RECT 23.18 415.53 695.02 417.24 ;
   RECT 23.18 417.24 695.02 418.95 ;
   RECT 23.18 418.95 695.02 420.66 ;
   RECT 23.18 420.66 695.02 422.37 ;
   RECT 23.18 422.37 695.02 424.08 ;
   RECT 23.18 424.08 695.02 425.79 ;
   RECT 23.18 425.79 695.02 427.5 ;
   RECT 23.18 427.5 695.02 429.21 ;
   RECT 23.18 429.21 695.02 430.92 ;
   RECT 23.18 430.92 695.02 432.63 ;
   RECT 23.18 432.63 695.02 434.34 ;
   RECT 23.18 434.34 695.02 436.05 ;
   RECT 23.18 436.05 695.02 437.76 ;
   RECT 23.18 437.76 695.02 439.47 ;
   RECT 23.18 439.47 695.02 441.18 ;
   RECT 23.18 441.18 695.02 442.89 ;
   RECT 23.18 442.89 695.02 444.6 ;
   RECT 23.18 444.6 695.02 446.31 ;
   RECT 23.18 446.31 695.02 448.02 ;
   RECT 23.18 448.02 695.02 449.73 ;
   RECT 23.18 449.73 695.02 451.44 ;
   RECT 23.18 451.44 695.02 453.15 ;
   RECT 23.18 453.15 695.02 454.86 ;
   RECT 23.18 454.86 695.02 456.57 ;
   RECT 23.18 456.57 695.02 458.28 ;
   RECT 23.18 458.28 695.02 459.99 ;
   RECT 23.18 459.99 695.02 461.7 ;
   RECT 23.18 461.7 695.02 463.41 ;
   RECT 23.18 463.41 695.02 465.12 ;
   RECT 23.18 465.12 695.02 466.83 ;
   RECT 23.18 466.83 695.02 468.54 ;
   RECT 23.18 468.54 695.02 470.25 ;
   RECT 23.18 470.25 695.02 471.96 ;
   RECT 23.18 471.96 695.02 473.67 ;
   RECT 23.18 473.67 695.02 475.38 ;
  LAYER via1 ;
   RECT 23.18 0.0 695.02 1.71 ;
   RECT 23.18 1.71 695.02 3.42 ;
   RECT 23.18 3.42 695.02 5.13 ;
   RECT 23.18 5.13 695.02 6.84 ;
   RECT 23.18 6.84 695.02 8.55 ;
   RECT 23.18 8.55 695.02 10.26 ;
   RECT 23.18 10.26 695.02 11.97 ;
   RECT 23.18 11.97 695.02 13.68 ;
   RECT 23.18 13.68 695.02 15.39 ;
   RECT 23.18 15.39 695.02 17.1 ;
   RECT 23.18 17.1 695.02 18.81 ;
   RECT 23.18 18.81 695.02 20.52 ;
   RECT 23.18 20.52 695.02 22.23 ;
   RECT 23.18 22.23 695.02 23.94 ;
   RECT 23.18 23.94 695.02 25.65 ;
   RECT 23.18 25.65 695.02 27.36 ;
   RECT 23.18 27.36 695.02 29.07 ;
   RECT 23.18 29.07 695.02 30.78 ;
   RECT 23.18 30.78 695.02 32.49 ;
   RECT 23.18 32.49 695.02 34.2 ;
   RECT 23.18 34.2 695.02 35.91 ;
   RECT 23.18 35.91 695.02 37.62 ;
   RECT 23.18 37.62 695.02 39.33 ;
   RECT 23.18 39.33 695.02 41.04 ;
   RECT 23.18 41.04 695.02 42.75 ;
   RECT 23.18 42.75 695.02 44.46 ;
   RECT 23.18 44.46 695.02 46.17 ;
   RECT 23.18 46.17 695.02 47.88 ;
   RECT 23.18 47.88 695.02 49.59 ;
   RECT 23.18 49.59 695.02 51.3 ;
   RECT 23.18 51.3 695.02 53.01 ;
   RECT 23.18 53.01 695.02 54.72 ;
   RECT 23.18 54.72 695.02 56.43 ;
   RECT 23.18 56.43 695.02 58.14 ;
   RECT 23.18 58.14 695.02 59.85 ;
   RECT 23.18 59.85 695.02 61.56 ;
   RECT 23.18 61.56 695.02 63.27 ;
   RECT 23.18 63.27 695.02 64.98 ;
   RECT 23.18 64.98 695.02 66.69 ;
   RECT 23.18 66.69 695.02 68.4 ;
   RECT 23.18 68.4 695.02 70.11 ;
   RECT 23.18 70.11 695.02 71.82 ;
   RECT 23.18 71.82 695.02 73.53 ;
   RECT 23.18 73.53 695.02 75.24 ;
   RECT 23.18 75.24 695.02 76.95 ;
   RECT 23.18 76.95 695.02 78.66 ;
   RECT 23.18 78.66 695.02 80.37 ;
   RECT 23.18 80.37 695.02 82.08 ;
   RECT 23.18 82.08 695.02 83.79 ;
   RECT 23.18 83.79 695.02 85.5 ;
   RECT 23.18 85.5 695.02 87.21 ;
   RECT 23.18 87.21 695.02 88.92 ;
   RECT 23.18 88.92 695.02 90.63 ;
   RECT 23.18 90.63 695.02 92.34 ;
   RECT 23.18 92.34 695.02 94.05 ;
   RECT 23.18 94.05 695.02 95.76 ;
   RECT 23.18 95.76 695.02 97.47 ;
   RECT 23.18 97.47 695.02 99.18 ;
   RECT 23.18 99.18 695.02 100.89 ;
   RECT 23.18 100.89 695.02 102.6 ;
   RECT 23.18 102.6 695.02 104.31 ;
   RECT 23.18 104.31 695.02 106.02 ;
   RECT 23.18 106.02 695.02 107.73 ;
   RECT 23.18 107.73 695.02 109.44 ;
   RECT 23.18 109.44 695.02 111.15 ;
   RECT 23.18 111.15 695.02 112.86 ;
   RECT 23.18 112.86 695.02 114.57 ;
   RECT 23.18 114.57 695.02 116.28 ;
   RECT 23.18 116.28 695.02 117.99 ;
   RECT 23.18 117.99 695.02 119.7 ;
   RECT 23.18 119.7 695.02 121.41 ;
   RECT 23.18 121.41 695.02 123.12 ;
   RECT 23.18 123.12 695.02 124.83 ;
   RECT 23.18 124.83 695.02 126.54 ;
   RECT 23.18 126.54 695.02 128.25 ;
   RECT 23.18 128.25 695.02 129.96 ;
   RECT 23.18 129.96 695.02 131.67 ;
   RECT 23.18 131.67 695.02 133.38 ;
   RECT 23.18 133.38 695.02 135.09 ;
   RECT 23.18 135.09 695.02 136.8 ;
   RECT 23.18 136.8 695.02 138.51 ;
   RECT 23.18 138.51 695.02 140.22 ;
   RECT 23.18 140.22 695.02 141.93 ;
   RECT 23.18 141.93 695.02 143.64 ;
   RECT 23.18 143.64 695.02 145.35 ;
   RECT 23.18 145.35 695.02 147.06 ;
   RECT 23.18 147.06 695.02 148.77 ;
   RECT 23.18 148.77 695.02 150.48 ;
   RECT 23.18 150.48 695.02 152.19 ;
   RECT 23.18 152.19 695.02 153.9 ;
   RECT 23.18 153.9 695.02 155.61 ;
   RECT 23.18 155.61 695.02 157.32 ;
   RECT 23.18 157.32 695.02 159.03 ;
   RECT 23.18 159.03 695.02 160.74 ;
   RECT 23.18 160.74 695.02 162.45 ;
   RECT 23.18 162.45 695.02 164.16 ;
   RECT 23.18 164.16 695.02 165.87 ;
   RECT 23.18 165.87 695.02 167.58 ;
   RECT 23.18 167.58 695.02 169.29 ;
   RECT 23.18 169.29 695.02 171.0 ;
   RECT 23.18 171.0 695.02 172.71 ;
   RECT 23.18 172.71 695.02 174.42 ;
   RECT 23.18 174.42 695.02 176.13 ;
   RECT 23.18 176.13 695.02 177.84 ;
   RECT 23.18 177.84 695.02 179.55 ;
   RECT 23.18 179.55 695.02 181.26 ;
   RECT 23.18 181.26 695.02 182.97 ;
   RECT 23.18 182.97 695.02 184.68 ;
   RECT 23.18 184.68 695.02 186.39 ;
   RECT 23.18 186.39 695.02 188.1 ;
   RECT 23.18 188.1 695.02 189.81 ;
   RECT 23.18 189.81 695.02 191.52 ;
   RECT 23.18 191.52 695.02 193.23 ;
   RECT 23.18 193.23 695.02 194.94 ;
   RECT 23.18 194.94 695.02 196.65 ;
   RECT 23.18 196.65 695.02 198.36 ;
   RECT 23.18 198.36 695.02 200.07 ;
   RECT 23.18 200.07 695.02 201.78 ;
   RECT 23.18 201.78 695.02 203.49 ;
   RECT 23.18 203.49 695.02 205.2 ;
   RECT 23.18 205.2 695.02 206.91 ;
   RECT 23.18 206.91 695.02 208.62 ;
   RECT 23.18 208.62 695.02 210.33 ;
   RECT 23.18 210.33 695.02 212.04 ;
   RECT 23.18 212.04 695.02 213.75 ;
   RECT 23.18 213.75 695.02 215.46 ;
   RECT 0.0 215.46 695.02 217.17 ;
   RECT 0.0 217.17 695.02 218.88 ;
   RECT 0.0 218.88 695.02 220.59 ;
   RECT 0.0 220.59 695.02 222.3 ;
   RECT 0.0 222.3 695.02 224.01 ;
   RECT 0.0 224.01 695.02 225.72 ;
   RECT 0.0 225.72 695.02 227.43 ;
   RECT 0.0 227.43 695.02 229.14 ;
   RECT 0.0 229.14 695.02 230.85 ;
   RECT 0.0 230.85 695.02 232.56 ;
   RECT 0.0 232.56 695.02 234.27 ;
   RECT 0.0 234.27 695.02 235.98 ;
   RECT 0.0 235.98 695.02 237.69 ;
   RECT 0.0 237.69 695.02 239.4 ;
   RECT 0.0 239.4 695.02 241.11 ;
   RECT 0.0 241.11 695.02 242.82 ;
   RECT 0.0 242.82 695.02 244.53 ;
   RECT 23.18 244.53 695.02 246.24 ;
   RECT 23.18 246.24 695.02 247.95 ;
   RECT 23.18 247.95 695.02 249.66 ;
   RECT 23.18 249.66 695.02 251.37 ;
   RECT 23.18 251.37 695.02 253.08 ;
   RECT 23.18 253.08 695.02 254.79 ;
   RECT 23.18 254.79 695.02 256.5 ;
   RECT 23.18 256.5 695.02 258.21 ;
   RECT 23.18 258.21 695.02 259.92 ;
   RECT 23.18 259.92 695.02 261.63 ;
   RECT 23.18 261.63 695.02 263.34 ;
   RECT 23.18 263.34 695.02 265.05 ;
   RECT 23.18 265.05 695.02 266.76 ;
   RECT 23.18 266.76 695.02 268.47 ;
   RECT 23.18 268.47 695.02 270.18 ;
   RECT 23.18 270.18 695.02 271.89 ;
   RECT 23.18 271.89 695.02 273.6 ;
   RECT 23.18 273.6 695.02 275.31 ;
   RECT 23.18 275.31 695.02 277.02 ;
   RECT 23.18 277.02 695.02 278.73 ;
   RECT 23.18 278.73 695.02 280.44 ;
   RECT 23.18 280.44 695.02 282.15 ;
   RECT 23.18 282.15 695.02 283.86 ;
   RECT 23.18 283.86 695.02 285.57 ;
   RECT 23.18 285.57 695.02 287.28 ;
   RECT 23.18 287.28 695.02 288.99 ;
   RECT 23.18 288.99 695.02 290.7 ;
   RECT 23.18 290.7 695.02 292.41 ;
   RECT 23.18 292.41 695.02 294.12 ;
   RECT 23.18 294.12 695.02 295.83 ;
   RECT 23.18 295.83 695.02 297.54 ;
   RECT 23.18 297.54 695.02 299.25 ;
   RECT 23.18 299.25 695.02 300.96 ;
   RECT 23.18 300.96 695.02 302.67 ;
   RECT 23.18 302.67 695.02 304.38 ;
   RECT 23.18 304.38 695.02 306.09 ;
   RECT 23.18 306.09 695.02 307.8 ;
   RECT 23.18 307.8 695.02 309.51 ;
   RECT 23.18 309.51 695.02 311.22 ;
   RECT 23.18 311.22 695.02 312.93 ;
   RECT 23.18 312.93 695.02 314.64 ;
   RECT 23.18 314.64 695.02 316.35 ;
   RECT 23.18 316.35 695.02 318.06 ;
   RECT 23.18 318.06 695.02 319.77 ;
   RECT 23.18 319.77 695.02 321.48 ;
   RECT 23.18 321.48 695.02 323.19 ;
   RECT 23.18 323.19 695.02 324.9 ;
   RECT 23.18 324.9 695.02 326.61 ;
   RECT 23.18 326.61 695.02 328.32 ;
   RECT 23.18 328.32 695.02 330.03 ;
   RECT 23.18 330.03 695.02 331.74 ;
   RECT 23.18 331.74 695.02 333.45 ;
   RECT 23.18 333.45 695.02 335.16 ;
   RECT 23.18 335.16 695.02 336.87 ;
   RECT 23.18 336.87 695.02 338.58 ;
   RECT 23.18 338.58 695.02 340.29 ;
   RECT 23.18 340.29 695.02 342.0 ;
   RECT 23.18 342.0 695.02 343.71 ;
   RECT 23.18 343.71 695.02 345.42 ;
   RECT 23.18 345.42 695.02 347.13 ;
   RECT 23.18 347.13 695.02 348.84 ;
   RECT 23.18 348.84 695.02 350.55 ;
   RECT 23.18 350.55 695.02 352.26 ;
   RECT 23.18 352.26 695.02 353.97 ;
   RECT 23.18 353.97 695.02 355.68 ;
   RECT 23.18 355.68 695.02 357.39 ;
   RECT 23.18 357.39 695.02 359.1 ;
   RECT 23.18 359.1 695.02 360.81 ;
   RECT 23.18 360.81 695.02 362.52 ;
   RECT 23.18 362.52 695.02 364.23 ;
   RECT 23.18 364.23 695.02 365.94 ;
   RECT 23.18 365.94 695.02 367.65 ;
   RECT 23.18 367.65 695.02 369.36 ;
   RECT 23.18 369.36 695.02 371.07 ;
   RECT 23.18 371.07 695.02 372.78 ;
   RECT 23.18 372.78 695.02 374.49 ;
   RECT 23.18 374.49 695.02 376.2 ;
   RECT 23.18 376.2 695.02 377.91 ;
   RECT 23.18 377.91 695.02 379.62 ;
   RECT 23.18 379.62 695.02 381.33 ;
   RECT 23.18 381.33 695.02 383.04 ;
   RECT 23.18 383.04 695.02 384.75 ;
   RECT 23.18 384.75 695.02 386.46 ;
   RECT 23.18 386.46 695.02 388.17 ;
   RECT 23.18 388.17 695.02 389.88 ;
   RECT 23.18 389.88 695.02 391.59 ;
   RECT 23.18 391.59 695.02 393.3 ;
   RECT 23.18 393.3 695.02 395.01 ;
   RECT 23.18 395.01 695.02 396.72 ;
   RECT 23.18 396.72 695.02 398.43 ;
   RECT 23.18 398.43 695.02 400.14 ;
   RECT 23.18 400.14 695.02 401.85 ;
   RECT 23.18 401.85 695.02 403.56 ;
   RECT 23.18 403.56 695.02 405.27 ;
   RECT 23.18 405.27 695.02 406.98 ;
   RECT 23.18 406.98 695.02 408.69 ;
   RECT 23.18 408.69 695.02 410.4 ;
   RECT 23.18 410.4 695.02 412.11 ;
   RECT 23.18 412.11 695.02 413.82 ;
   RECT 23.18 413.82 695.02 415.53 ;
   RECT 23.18 415.53 695.02 417.24 ;
   RECT 23.18 417.24 695.02 418.95 ;
   RECT 23.18 418.95 695.02 420.66 ;
   RECT 23.18 420.66 695.02 422.37 ;
   RECT 23.18 422.37 695.02 424.08 ;
   RECT 23.18 424.08 695.02 425.79 ;
   RECT 23.18 425.79 695.02 427.5 ;
   RECT 23.18 427.5 695.02 429.21 ;
   RECT 23.18 429.21 695.02 430.92 ;
   RECT 23.18 430.92 695.02 432.63 ;
   RECT 23.18 432.63 695.02 434.34 ;
   RECT 23.18 434.34 695.02 436.05 ;
   RECT 23.18 436.05 695.02 437.76 ;
   RECT 23.18 437.76 695.02 439.47 ;
   RECT 23.18 439.47 695.02 441.18 ;
   RECT 23.18 441.18 695.02 442.89 ;
   RECT 23.18 442.89 695.02 444.6 ;
   RECT 23.18 444.6 695.02 446.31 ;
   RECT 23.18 446.31 695.02 448.02 ;
   RECT 23.18 448.02 695.02 449.73 ;
   RECT 23.18 449.73 695.02 451.44 ;
   RECT 23.18 451.44 695.02 453.15 ;
   RECT 23.18 453.15 695.02 454.86 ;
   RECT 23.18 454.86 695.02 456.57 ;
   RECT 23.18 456.57 695.02 458.28 ;
   RECT 23.18 458.28 695.02 459.99 ;
   RECT 23.18 459.99 695.02 461.7 ;
   RECT 23.18 461.7 695.02 463.41 ;
   RECT 23.18 463.41 695.02 465.12 ;
   RECT 23.18 465.12 695.02 466.83 ;
   RECT 23.18 466.83 695.02 468.54 ;
   RECT 23.18 468.54 695.02 470.25 ;
   RECT 23.18 470.25 695.02 471.96 ;
   RECT 23.18 471.96 695.02 473.67 ;
   RECT 23.18 473.67 695.02 475.38 ;
  LAYER metal2 ;
   RECT 23.18 0.0 695.02 1.71 ;
   RECT 23.18 1.71 695.02 3.42 ;
   RECT 23.18 3.42 695.02 5.13 ;
   RECT 23.18 5.13 695.02 6.84 ;
   RECT 23.18 6.84 695.02 8.55 ;
   RECT 23.18 8.55 695.02 10.26 ;
   RECT 23.18 10.26 695.02 11.97 ;
   RECT 23.18 11.97 695.02 13.68 ;
   RECT 23.18 13.68 695.02 15.39 ;
   RECT 23.18 15.39 695.02 17.1 ;
   RECT 23.18 17.1 695.02 18.81 ;
   RECT 23.18 18.81 695.02 20.52 ;
   RECT 23.18 20.52 695.02 22.23 ;
   RECT 23.18 22.23 695.02 23.94 ;
   RECT 23.18 23.94 695.02 25.65 ;
   RECT 23.18 25.65 695.02 27.36 ;
   RECT 23.18 27.36 695.02 29.07 ;
   RECT 23.18 29.07 695.02 30.78 ;
   RECT 23.18 30.78 695.02 32.49 ;
   RECT 23.18 32.49 695.02 34.2 ;
   RECT 23.18 34.2 695.02 35.91 ;
   RECT 23.18 35.91 695.02 37.62 ;
   RECT 23.18 37.62 695.02 39.33 ;
   RECT 23.18 39.33 695.02 41.04 ;
   RECT 23.18 41.04 695.02 42.75 ;
   RECT 23.18 42.75 695.02 44.46 ;
   RECT 23.18 44.46 695.02 46.17 ;
   RECT 23.18 46.17 695.02 47.88 ;
   RECT 23.18 47.88 695.02 49.59 ;
   RECT 23.18 49.59 695.02 51.3 ;
   RECT 23.18 51.3 695.02 53.01 ;
   RECT 23.18 53.01 695.02 54.72 ;
   RECT 23.18 54.72 695.02 56.43 ;
   RECT 23.18 56.43 695.02 58.14 ;
   RECT 23.18 58.14 695.02 59.85 ;
   RECT 23.18 59.85 695.02 61.56 ;
   RECT 23.18 61.56 695.02 63.27 ;
   RECT 23.18 63.27 695.02 64.98 ;
   RECT 23.18 64.98 695.02 66.69 ;
   RECT 23.18 66.69 695.02 68.4 ;
   RECT 23.18 68.4 695.02 70.11 ;
   RECT 23.18 70.11 695.02 71.82 ;
   RECT 23.18 71.82 695.02 73.53 ;
   RECT 23.18 73.53 695.02 75.24 ;
   RECT 23.18 75.24 695.02 76.95 ;
   RECT 23.18 76.95 695.02 78.66 ;
   RECT 23.18 78.66 695.02 80.37 ;
   RECT 23.18 80.37 695.02 82.08 ;
   RECT 23.18 82.08 695.02 83.79 ;
   RECT 23.18 83.79 695.02 85.5 ;
   RECT 23.18 85.5 695.02 87.21 ;
   RECT 23.18 87.21 695.02 88.92 ;
   RECT 23.18 88.92 695.02 90.63 ;
   RECT 23.18 90.63 695.02 92.34 ;
   RECT 23.18 92.34 695.02 94.05 ;
   RECT 23.18 94.05 695.02 95.76 ;
   RECT 23.18 95.76 695.02 97.47 ;
   RECT 23.18 97.47 695.02 99.18 ;
   RECT 23.18 99.18 695.02 100.89 ;
   RECT 23.18 100.89 695.02 102.6 ;
   RECT 23.18 102.6 695.02 104.31 ;
   RECT 23.18 104.31 695.02 106.02 ;
   RECT 23.18 106.02 695.02 107.73 ;
   RECT 23.18 107.73 695.02 109.44 ;
   RECT 23.18 109.44 695.02 111.15 ;
   RECT 23.18 111.15 695.02 112.86 ;
   RECT 23.18 112.86 695.02 114.57 ;
   RECT 23.18 114.57 695.02 116.28 ;
   RECT 23.18 116.28 695.02 117.99 ;
   RECT 23.18 117.99 695.02 119.7 ;
   RECT 23.18 119.7 695.02 121.41 ;
   RECT 23.18 121.41 695.02 123.12 ;
   RECT 23.18 123.12 695.02 124.83 ;
   RECT 23.18 124.83 695.02 126.54 ;
   RECT 23.18 126.54 695.02 128.25 ;
   RECT 23.18 128.25 695.02 129.96 ;
   RECT 23.18 129.96 695.02 131.67 ;
   RECT 23.18 131.67 695.02 133.38 ;
   RECT 23.18 133.38 695.02 135.09 ;
   RECT 23.18 135.09 695.02 136.8 ;
   RECT 23.18 136.8 695.02 138.51 ;
   RECT 23.18 138.51 695.02 140.22 ;
   RECT 23.18 140.22 695.02 141.93 ;
   RECT 23.18 141.93 695.02 143.64 ;
   RECT 23.18 143.64 695.02 145.35 ;
   RECT 23.18 145.35 695.02 147.06 ;
   RECT 23.18 147.06 695.02 148.77 ;
   RECT 23.18 148.77 695.02 150.48 ;
   RECT 23.18 150.48 695.02 152.19 ;
   RECT 23.18 152.19 695.02 153.9 ;
   RECT 23.18 153.9 695.02 155.61 ;
   RECT 23.18 155.61 695.02 157.32 ;
   RECT 23.18 157.32 695.02 159.03 ;
   RECT 23.18 159.03 695.02 160.74 ;
   RECT 23.18 160.74 695.02 162.45 ;
   RECT 23.18 162.45 695.02 164.16 ;
   RECT 23.18 164.16 695.02 165.87 ;
   RECT 23.18 165.87 695.02 167.58 ;
   RECT 23.18 167.58 695.02 169.29 ;
   RECT 23.18 169.29 695.02 171.0 ;
   RECT 23.18 171.0 695.02 172.71 ;
   RECT 23.18 172.71 695.02 174.42 ;
   RECT 23.18 174.42 695.02 176.13 ;
   RECT 23.18 176.13 695.02 177.84 ;
   RECT 23.18 177.84 695.02 179.55 ;
   RECT 23.18 179.55 695.02 181.26 ;
   RECT 23.18 181.26 695.02 182.97 ;
   RECT 23.18 182.97 695.02 184.68 ;
   RECT 23.18 184.68 695.02 186.39 ;
   RECT 23.18 186.39 695.02 188.1 ;
   RECT 23.18 188.1 695.02 189.81 ;
   RECT 23.18 189.81 695.02 191.52 ;
   RECT 23.18 191.52 695.02 193.23 ;
   RECT 23.18 193.23 695.02 194.94 ;
   RECT 23.18 194.94 695.02 196.65 ;
   RECT 23.18 196.65 695.02 198.36 ;
   RECT 23.18 198.36 695.02 200.07 ;
   RECT 23.18 200.07 695.02 201.78 ;
   RECT 23.18 201.78 695.02 203.49 ;
   RECT 23.18 203.49 695.02 205.2 ;
   RECT 23.18 205.2 695.02 206.91 ;
   RECT 23.18 206.91 695.02 208.62 ;
   RECT 23.18 208.62 695.02 210.33 ;
   RECT 23.18 210.33 695.02 212.04 ;
   RECT 23.18 212.04 695.02 213.75 ;
   RECT 23.18 213.75 695.02 215.46 ;
   RECT 0.0 215.46 695.02 217.17 ;
   RECT 0.0 217.17 695.02 218.88 ;
   RECT 0.0 218.88 695.02 220.59 ;
   RECT 0.0 220.59 695.02 222.3 ;
   RECT 0.0 222.3 695.02 224.01 ;
   RECT 0.0 224.01 695.02 225.72 ;
   RECT 0.0 225.72 695.02 227.43 ;
   RECT 0.0 227.43 695.02 229.14 ;
   RECT 0.0 229.14 695.02 230.85 ;
   RECT 0.0 230.85 695.02 232.56 ;
   RECT 0.0 232.56 695.02 234.27 ;
   RECT 0.0 234.27 695.02 235.98 ;
   RECT 0.0 235.98 695.02 237.69 ;
   RECT 0.0 237.69 695.02 239.4 ;
   RECT 0.0 239.4 695.02 241.11 ;
   RECT 0.0 241.11 695.02 242.82 ;
   RECT 0.0 242.82 695.02 244.53 ;
   RECT 23.18 244.53 695.02 246.24 ;
   RECT 23.18 246.24 695.02 247.95 ;
   RECT 23.18 247.95 695.02 249.66 ;
   RECT 23.18 249.66 695.02 251.37 ;
   RECT 23.18 251.37 695.02 253.08 ;
   RECT 23.18 253.08 695.02 254.79 ;
   RECT 23.18 254.79 695.02 256.5 ;
   RECT 23.18 256.5 695.02 258.21 ;
   RECT 23.18 258.21 695.02 259.92 ;
   RECT 23.18 259.92 695.02 261.63 ;
   RECT 23.18 261.63 695.02 263.34 ;
   RECT 23.18 263.34 695.02 265.05 ;
   RECT 23.18 265.05 695.02 266.76 ;
   RECT 23.18 266.76 695.02 268.47 ;
   RECT 23.18 268.47 695.02 270.18 ;
   RECT 23.18 270.18 695.02 271.89 ;
   RECT 23.18 271.89 695.02 273.6 ;
   RECT 23.18 273.6 695.02 275.31 ;
   RECT 23.18 275.31 695.02 277.02 ;
   RECT 23.18 277.02 695.02 278.73 ;
   RECT 23.18 278.73 695.02 280.44 ;
   RECT 23.18 280.44 695.02 282.15 ;
   RECT 23.18 282.15 695.02 283.86 ;
   RECT 23.18 283.86 695.02 285.57 ;
   RECT 23.18 285.57 695.02 287.28 ;
   RECT 23.18 287.28 695.02 288.99 ;
   RECT 23.18 288.99 695.02 290.7 ;
   RECT 23.18 290.7 695.02 292.41 ;
   RECT 23.18 292.41 695.02 294.12 ;
   RECT 23.18 294.12 695.02 295.83 ;
   RECT 23.18 295.83 695.02 297.54 ;
   RECT 23.18 297.54 695.02 299.25 ;
   RECT 23.18 299.25 695.02 300.96 ;
   RECT 23.18 300.96 695.02 302.67 ;
   RECT 23.18 302.67 695.02 304.38 ;
   RECT 23.18 304.38 695.02 306.09 ;
   RECT 23.18 306.09 695.02 307.8 ;
   RECT 23.18 307.8 695.02 309.51 ;
   RECT 23.18 309.51 695.02 311.22 ;
   RECT 23.18 311.22 695.02 312.93 ;
   RECT 23.18 312.93 695.02 314.64 ;
   RECT 23.18 314.64 695.02 316.35 ;
   RECT 23.18 316.35 695.02 318.06 ;
   RECT 23.18 318.06 695.02 319.77 ;
   RECT 23.18 319.77 695.02 321.48 ;
   RECT 23.18 321.48 695.02 323.19 ;
   RECT 23.18 323.19 695.02 324.9 ;
   RECT 23.18 324.9 695.02 326.61 ;
   RECT 23.18 326.61 695.02 328.32 ;
   RECT 23.18 328.32 695.02 330.03 ;
   RECT 23.18 330.03 695.02 331.74 ;
   RECT 23.18 331.74 695.02 333.45 ;
   RECT 23.18 333.45 695.02 335.16 ;
   RECT 23.18 335.16 695.02 336.87 ;
   RECT 23.18 336.87 695.02 338.58 ;
   RECT 23.18 338.58 695.02 340.29 ;
   RECT 23.18 340.29 695.02 342.0 ;
   RECT 23.18 342.0 695.02 343.71 ;
   RECT 23.18 343.71 695.02 345.42 ;
   RECT 23.18 345.42 695.02 347.13 ;
   RECT 23.18 347.13 695.02 348.84 ;
   RECT 23.18 348.84 695.02 350.55 ;
   RECT 23.18 350.55 695.02 352.26 ;
   RECT 23.18 352.26 695.02 353.97 ;
   RECT 23.18 353.97 695.02 355.68 ;
   RECT 23.18 355.68 695.02 357.39 ;
   RECT 23.18 357.39 695.02 359.1 ;
   RECT 23.18 359.1 695.02 360.81 ;
   RECT 23.18 360.81 695.02 362.52 ;
   RECT 23.18 362.52 695.02 364.23 ;
   RECT 23.18 364.23 695.02 365.94 ;
   RECT 23.18 365.94 695.02 367.65 ;
   RECT 23.18 367.65 695.02 369.36 ;
   RECT 23.18 369.36 695.02 371.07 ;
   RECT 23.18 371.07 695.02 372.78 ;
   RECT 23.18 372.78 695.02 374.49 ;
   RECT 23.18 374.49 695.02 376.2 ;
   RECT 23.18 376.2 695.02 377.91 ;
   RECT 23.18 377.91 695.02 379.62 ;
   RECT 23.18 379.62 695.02 381.33 ;
   RECT 23.18 381.33 695.02 383.04 ;
   RECT 23.18 383.04 695.02 384.75 ;
   RECT 23.18 384.75 695.02 386.46 ;
   RECT 23.18 386.46 695.02 388.17 ;
   RECT 23.18 388.17 695.02 389.88 ;
   RECT 23.18 389.88 695.02 391.59 ;
   RECT 23.18 391.59 695.02 393.3 ;
   RECT 23.18 393.3 695.02 395.01 ;
   RECT 23.18 395.01 695.02 396.72 ;
   RECT 23.18 396.72 695.02 398.43 ;
   RECT 23.18 398.43 695.02 400.14 ;
   RECT 23.18 400.14 695.02 401.85 ;
   RECT 23.18 401.85 695.02 403.56 ;
   RECT 23.18 403.56 695.02 405.27 ;
   RECT 23.18 405.27 695.02 406.98 ;
   RECT 23.18 406.98 695.02 408.69 ;
   RECT 23.18 408.69 695.02 410.4 ;
   RECT 23.18 410.4 695.02 412.11 ;
   RECT 23.18 412.11 695.02 413.82 ;
   RECT 23.18 413.82 695.02 415.53 ;
   RECT 23.18 415.53 695.02 417.24 ;
   RECT 23.18 417.24 695.02 418.95 ;
   RECT 23.18 418.95 695.02 420.66 ;
   RECT 23.18 420.66 695.02 422.37 ;
   RECT 23.18 422.37 695.02 424.08 ;
   RECT 23.18 424.08 695.02 425.79 ;
   RECT 23.18 425.79 695.02 427.5 ;
   RECT 23.18 427.5 695.02 429.21 ;
   RECT 23.18 429.21 695.02 430.92 ;
   RECT 23.18 430.92 695.02 432.63 ;
   RECT 23.18 432.63 695.02 434.34 ;
   RECT 23.18 434.34 695.02 436.05 ;
   RECT 23.18 436.05 695.02 437.76 ;
   RECT 23.18 437.76 695.02 439.47 ;
   RECT 23.18 439.47 695.02 441.18 ;
   RECT 23.18 441.18 695.02 442.89 ;
   RECT 23.18 442.89 695.02 444.6 ;
   RECT 23.18 444.6 695.02 446.31 ;
   RECT 23.18 446.31 695.02 448.02 ;
   RECT 23.18 448.02 695.02 449.73 ;
   RECT 23.18 449.73 695.02 451.44 ;
   RECT 23.18 451.44 695.02 453.15 ;
   RECT 23.18 453.15 695.02 454.86 ;
   RECT 23.18 454.86 695.02 456.57 ;
   RECT 23.18 456.57 695.02 458.28 ;
   RECT 23.18 458.28 695.02 459.99 ;
   RECT 23.18 459.99 695.02 461.7 ;
   RECT 23.18 461.7 695.02 463.41 ;
   RECT 23.18 463.41 695.02 465.12 ;
   RECT 23.18 465.12 695.02 466.83 ;
   RECT 23.18 466.83 695.02 468.54 ;
   RECT 23.18 468.54 695.02 470.25 ;
   RECT 23.18 470.25 695.02 471.96 ;
   RECT 23.18 471.96 695.02 473.67 ;
   RECT 23.18 473.67 695.02 475.38 ;
  LAYER via2 ;
   RECT 23.18 0.0 695.02 1.71 ;
   RECT 23.18 1.71 695.02 3.42 ;
   RECT 23.18 3.42 695.02 5.13 ;
   RECT 23.18 5.13 695.02 6.84 ;
   RECT 23.18 6.84 695.02 8.55 ;
   RECT 23.18 8.55 695.02 10.26 ;
   RECT 23.18 10.26 695.02 11.97 ;
   RECT 23.18 11.97 695.02 13.68 ;
   RECT 23.18 13.68 695.02 15.39 ;
   RECT 23.18 15.39 695.02 17.1 ;
   RECT 23.18 17.1 695.02 18.81 ;
   RECT 23.18 18.81 695.02 20.52 ;
   RECT 23.18 20.52 695.02 22.23 ;
   RECT 23.18 22.23 695.02 23.94 ;
   RECT 23.18 23.94 695.02 25.65 ;
   RECT 23.18 25.65 695.02 27.36 ;
   RECT 23.18 27.36 695.02 29.07 ;
   RECT 23.18 29.07 695.02 30.78 ;
   RECT 23.18 30.78 695.02 32.49 ;
   RECT 23.18 32.49 695.02 34.2 ;
   RECT 23.18 34.2 695.02 35.91 ;
   RECT 23.18 35.91 695.02 37.62 ;
   RECT 23.18 37.62 695.02 39.33 ;
   RECT 23.18 39.33 695.02 41.04 ;
   RECT 23.18 41.04 695.02 42.75 ;
   RECT 23.18 42.75 695.02 44.46 ;
   RECT 23.18 44.46 695.02 46.17 ;
   RECT 23.18 46.17 695.02 47.88 ;
   RECT 23.18 47.88 695.02 49.59 ;
   RECT 23.18 49.59 695.02 51.3 ;
   RECT 23.18 51.3 695.02 53.01 ;
   RECT 23.18 53.01 695.02 54.72 ;
   RECT 23.18 54.72 695.02 56.43 ;
   RECT 23.18 56.43 695.02 58.14 ;
   RECT 23.18 58.14 695.02 59.85 ;
   RECT 23.18 59.85 695.02 61.56 ;
   RECT 23.18 61.56 695.02 63.27 ;
   RECT 23.18 63.27 695.02 64.98 ;
   RECT 23.18 64.98 695.02 66.69 ;
   RECT 23.18 66.69 695.02 68.4 ;
   RECT 23.18 68.4 695.02 70.11 ;
   RECT 23.18 70.11 695.02 71.82 ;
   RECT 23.18 71.82 695.02 73.53 ;
   RECT 23.18 73.53 695.02 75.24 ;
   RECT 23.18 75.24 695.02 76.95 ;
   RECT 23.18 76.95 695.02 78.66 ;
   RECT 23.18 78.66 695.02 80.37 ;
   RECT 23.18 80.37 695.02 82.08 ;
   RECT 23.18 82.08 695.02 83.79 ;
   RECT 23.18 83.79 695.02 85.5 ;
   RECT 23.18 85.5 695.02 87.21 ;
   RECT 23.18 87.21 695.02 88.92 ;
   RECT 23.18 88.92 695.02 90.63 ;
   RECT 23.18 90.63 695.02 92.34 ;
   RECT 23.18 92.34 695.02 94.05 ;
   RECT 23.18 94.05 695.02 95.76 ;
   RECT 23.18 95.76 695.02 97.47 ;
   RECT 23.18 97.47 695.02 99.18 ;
   RECT 23.18 99.18 695.02 100.89 ;
   RECT 23.18 100.89 695.02 102.6 ;
   RECT 23.18 102.6 695.02 104.31 ;
   RECT 23.18 104.31 695.02 106.02 ;
   RECT 23.18 106.02 695.02 107.73 ;
   RECT 23.18 107.73 695.02 109.44 ;
   RECT 23.18 109.44 695.02 111.15 ;
   RECT 23.18 111.15 695.02 112.86 ;
   RECT 23.18 112.86 695.02 114.57 ;
   RECT 23.18 114.57 695.02 116.28 ;
   RECT 23.18 116.28 695.02 117.99 ;
   RECT 23.18 117.99 695.02 119.7 ;
   RECT 23.18 119.7 695.02 121.41 ;
   RECT 23.18 121.41 695.02 123.12 ;
   RECT 23.18 123.12 695.02 124.83 ;
   RECT 23.18 124.83 695.02 126.54 ;
   RECT 23.18 126.54 695.02 128.25 ;
   RECT 23.18 128.25 695.02 129.96 ;
   RECT 23.18 129.96 695.02 131.67 ;
   RECT 23.18 131.67 695.02 133.38 ;
   RECT 23.18 133.38 695.02 135.09 ;
   RECT 23.18 135.09 695.02 136.8 ;
   RECT 23.18 136.8 695.02 138.51 ;
   RECT 23.18 138.51 695.02 140.22 ;
   RECT 23.18 140.22 695.02 141.93 ;
   RECT 23.18 141.93 695.02 143.64 ;
   RECT 23.18 143.64 695.02 145.35 ;
   RECT 23.18 145.35 695.02 147.06 ;
   RECT 23.18 147.06 695.02 148.77 ;
   RECT 23.18 148.77 695.02 150.48 ;
   RECT 23.18 150.48 695.02 152.19 ;
   RECT 23.18 152.19 695.02 153.9 ;
   RECT 23.18 153.9 695.02 155.61 ;
   RECT 23.18 155.61 695.02 157.32 ;
   RECT 23.18 157.32 695.02 159.03 ;
   RECT 23.18 159.03 695.02 160.74 ;
   RECT 23.18 160.74 695.02 162.45 ;
   RECT 23.18 162.45 695.02 164.16 ;
   RECT 23.18 164.16 695.02 165.87 ;
   RECT 23.18 165.87 695.02 167.58 ;
   RECT 23.18 167.58 695.02 169.29 ;
   RECT 23.18 169.29 695.02 171.0 ;
   RECT 23.18 171.0 695.02 172.71 ;
   RECT 23.18 172.71 695.02 174.42 ;
   RECT 23.18 174.42 695.02 176.13 ;
   RECT 23.18 176.13 695.02 177.84 ;
   RECT 23.18 177.84 695.02 179.55 ;
   RECT 23.18 179.55 695.02 181.26 ;
   RECT 23.18 181.26 695.02 182.97 ;
   RECT 23.18 182.97 695.02 184.68 ;
   RECT 23.18 184.68 695.02 186.39 ;
   RECT 23.18 186.39 695.02 188.1 ;
   RECT 23.18 188.1 695.02 189.81 ;
   RECT 23.18 189.81 695.02 191.52 ;
   RECT 23.18 191.52 695.02 193.23 ;
   RECT 23.18 193.23 695.02 194.94 ;
   RECT 23.18 194.94 695.02 196.65 ;
   RECT 23.18 196.65 695.02 198.36 ;
   RECT 23.18 198.36 695.02 200.07 ;
   RECT 23.18 200.07 695.02 201.78 ;
   RECT 23.18 201.78 695.02 203.49 ;
   RECT 23.18 203.49 695.02 205.2 ;
   RECT 23.18 205.2 695.02 206.91 ;
   RECT 23.18 206.91 695.02 208.62 ;
   RECT 23.18 208.62 695.02 210.33 ;
   RECT 23.18 210.33 695.02 212.04 ;
   RECT 23.18 212.04 695.02 213.75 ;
   RECT 23.18 213.75 695.02 215.46 ;
   RECT 0.0 215.46 695.02 217.17 ;
   RECT 0.0 217.17 695.02 218.88 ;
   RECT 0.0 218.88 695.02 220.59 ;
   RECT 0.0 220.59 695.02 222.3 ;
   RECT 0.0 222.3 695.02 224.01 ;
   RECT 0.0 224.01 695.02 225.72 ;
   RECT 0.0 225.72 695.02 227.43 ;
   RECT 0.0 227.43 695.02 229.14 ;
   RECT 0.0 229.14 695.02 230.85 ;
   RECT 0.0 230.85 695.02 232.56 ;
   RECT 0.0 232.56 695.02 234.27 ;
   RECT 0.0 234.27 695.02 235.98 ;
   RECT 0.0 235.98 695.02 237.69 ;
   RECT 0.0 237.69 695.02 239.4 ;
   RECT 0.0 239.4 695.02 241.11 ;
   RECT 0.0 241.11 695.02 242.82 ;
   RECT 0.0 242.82 695.02 244.53 ;
   RECT 23.18 244.53 695.02 246.24 ;
   RECT 23.18 246.24 695.02 247.95 ;
   RECT 23.18 247.95 695.02 249.66 ;
   RECT 23.18 249.66 695.02 251.37 ;
   RECT 23.18 251.37 695.02 253.08 ;
   RECT 23.18 253.08 695.02 254.79 ;
   RECT 23.18 254.79 695.02 256.5 ;
   RECT 23.18 256.5 695.02 258.21 ;
   RECT 23.18 258.21 695.02 259.92 ;
   RECT 23.18 259.92 695.02 261.63 ;
   RECT 23.18 261.63 695.02 263.34 ;
   RECT 23.18 263.34 695.02 265.05 ;
   RECT 23.18 265.05 695.02 266.76 ;
   RECT 23.18 266.76 695.02 268.47 ;
   RECT 23.18 268.47 695.02 270.18 ;
   RECT 23.18 270.18 695.02 271.89 ;
   RECT 23.18 271.89 695.02 273.6 ;
   RECT 23.18 273.6 695.02 275.31 ;
   RECT 23.18 275.31 695.02 277.02 ;
   RECT 23.18 277.02 695.02 278.73 ;
   RECT 23.18 278.73 695.02 280.44 ;
   RECT 23.18 280.44 695.02 282.15 ;
   RECT 23.18 282.15 695.02 283.86 ;
   RECT 23.18 283.86 695.02 285.57 ;
   RECT 23.18 285.57 695.02 287.28 ;
   RECT 23.18 287.28 695.02 288.99 ;
   RECT 23.18 288.99 695.02 290.7 ;
   RECT 23.18 290.7 695.02 292.41 ;
   RECT 23.18 292.41 695.02 294.12 ;
   RECT 23.18 294.12 695.02 295.83 ;
   RECT 23.18 295.83 695.02 297.54 ;
   RECT 23.18 297.54 695.02 299.25 ;
   RECT 23.18 299.25 695.02 300.96 ;
   RECT 23.18 300.96 695.02 302.67 ;
   RECT 23.18 302.67 695.02 304.38 ;
   RECT 23.18 304.38 695.02 306.09 ;
   RECT 23.18 306.09 695.02 307.8 ;
   RECT 23.18 307.8 695.02 309.51 ;
   RECT 23.18 309.51 695.02 311.22 ;
   RECT 23.18 311.22 695.02 312.93 ;
   RECT 23.18 312.93 695.02 314.64 ;
   RECT 23.18 314.64 695.02 316.35 ;
   RECT 23.18 316.35 695.02 318.06 ;
   RECT 23.18 318.06 695.02 319.77 ;
   RECT 23.18 319.77 695.02 321.48 ;
   RECT 23.18 321.48 695.02 323.19 ;
   RECT 23.18 323.19 695.02 324.9 ;
   RECT 23.18 324.9 695.02 326.61 ;
   RECT 23.18 326.61 695.02 328.32 ;
   RECT 23.18 328.32 695.02 330.03 ;
   RECT 23.18 330.03 695.02 331.74 ;
   RECT 23.18 331.74 695.02 333.45 ;
   RECT 23.18 333.45 695.02 335.16 ;
   RECT 23.18 335.16 695.02 336.87 ;
   RECT 23.18 336.87 695.02 338.58 ;
   RECT 23.18 338.58 695.02 340.29 ;
   RECT 23.18 340.29 695.02 342.0 ;
   RECT 23.18 342.0 695.02 343.71 ;
   RECT 23.18 343.71 695.02 345.42 ;
   RECT 23.18 345.42 695.02 347.13 ;
   RECT 23.18 347.13 695.02 348.84 ;
   RECT 23.18 348.84 695.02 350.55 ;
   RECT 23.18 350.55 695.02 352.26 ;
   RECT 23.18 352.26 695.02 353.97 ;
   RECT 23.18 353.97 695.02 355.68 ;
   RECT 23.18 355.68 695.02 357.39 ;
   RECT 23.18 357.39 695.02 359.1 ;
   RECT 23.18 359.1 695.02 360.81 ;
   RECT 23.18 360.81 695.02 362.52 ;
   RECT 23.18 362.52 695.02 364.23 ;
   RECT 23.18 364.23 695.02 365.94 ;
   RECT 23.18 365.94 695.02 367.65 ;
   RECT 23.18 367.65 695.02 369.36 ;
   RECT 23.18 369.36 695.02 371.07 ;
   RECT 23.18 371.07 695.02 372.78 ;
   RECT 23.18 372.78 695.02 374.49 ;
   RECT 23.18 374.49 695.02 376.2 ;
   RECT 23.18 376.2 695.02 377.91 ;
   RECT 23.18 377.91 695.02 379.62 ;
   RECT 23.18 379.62 695.02 381.33 ;
   RECT 23.18 381.33 695.02 383.04 ;
   RECT 23.18 383.04 695.02 384.75 ;
   RECT 23.18 384.75 695.02 386.46 ;
   RECT 23.18 386.46 695.02 388.17 ;
   RECT 23.18 388.17 695.02 389.88 ;
   RECT 23.18 389.88 695.02 391.59 ;
   RECT 23.18 391.59 695.02 393.3 ;
   RECT 23.18 393.3 695.02 395.01 ;
   RECT 23.18 395.01 695.02 396.72 ;
   RECT 23.18 396.72 695.02 398.43 ;
   RECT 23.18 398.43 695.02 400.14 ;
   RECT 23.18 400.14 695.02 401.85 ;
   RECT 23.18 401.85 695.02 403.56 ;
   RECT 23.18 403.56 695.02 405.27 ;
   RECT 23.18 405.27 695.02 406.98 ;
   RECT 23.18 406.98 695.02 408.69 ;
   RECT 23.18 408.69 695.02 410.4 ;
   RECT 23.18 410.4 695.02 412.11 ;
   RECT 23.18 412.11 695.02 413.82 ;
   RECT 23.18 413.82 695.02 415.53 ;
   RECT 23.18 415.53 695.02 417.24 ;
   RECT 23.18 417.24 695.02 418.95 ;
   RECT 23.18 418.95 695.02 420.66 ;
   RECT 23.18 420.66 695.02 422.37 ;
   RECT 23.18 422.37 695.02 424.08 ;
   RECT 23.18 424.08 695.02 425.79 ;
   RECT 23.18 425.79 695.02 427.5 ;
   RECT 23.18 427.5 695.02 429.21 ;
   RECT 23.18 429.21 695.02 430.92 ;
   RECT 23.18 430.92 695.02 432.63 ;
   RECT 23.18 432.63 695.02 434.34 ;
   RECT 23.18 434.34 695.02 436.05 ;
   RECT 23.18 436.05 695.02 437.76 ;
   RECT 23.18 437.76 695.02 439.47 ;
   RECT 23.18 439.47 695.02 441.18 ;
   RECT 23.18 441.18 695.02 442.89 ;
   RECT 23.18 442.89 695.02 444.6 ;
   RECT 23.18 444.6 695.02 446.31 ;
   RECT 23.18 446.31 695.02 448.02 ;
   RECT 23.18 448.02 695.02 449.73 ;
   RECT 23.18 449.73 695.02 451.44 ;
   RECT 23.18 451.44 695.02 453.15 ;
   RECT 23.18 453.15 695.02 454.86 ;
   RECT 23.18 454.86 695.02 456.57 ;
   RECT 23.18 456.57 695.02 458.28 ;
   RECT 23.18 458.28 695.02 459.99 ;
   RECT 23.18 459.99 695.02 461.7 ;
   RECT 23.18 461.7 695.02 463.41 ;
   RECT 23.18 463.41 695.02 465.12 ;
   RECT 23.18 465.12 695.02 466.83 ;
   RECT 23.18 466.83 695.02 468.54 ;
   RECT 23.18 468.54 695.02 470.25 ;
   RECT 23.18 470.25 695.02 471.96 ;
   RECT 23.18 471.96 695.02 473.67 ;
   RECT 23.18 473.67 695.02 475.38 ;
  LAYER metal3 ;
   RECT 23.18 0.0 695.02 1.71 ;
   RECT 23.18 1.71 695.02 3.42 ;
   RECT 23.18 3.42 695.02 5.13 ;
   RECT 23.18 5.13 695.02 6.84 ;
   RECT 23.18 6.84 695.02 8.55 ;
   RECT 23.18 8.55 695.02 10.26 ;
   RECT 23.18 10.26 695.02 11.97 ;
   RECT 23.18 11.97 695.02 13.68 ;
   RECT 23.18 13.68 695.02 15.39 ;
   RECT 23.18 15.39 695.02 17.1 ;
   RECT 23.18 17.1 695.02 18.81 ;
   RECT 23.18 18.81 695.02 20.52 ;
   RECT 23.18 20.52 695.02 22.23 ;
   RECT 23.18 22.23 695.02 23.94 ;
   RECT 23.18 23.94 695.02 25.65 ;
   RECT 23.18 25.65 695.02 27.36 ;
   RECT 23.18 27.36 695.02 29.07 ;
   RECT 23.18 29.07 695.02 30.78 ;
   RECT 23.18 30.78 695.02 32.49 ;
   RECT 23.18 32.49 695.02 34.2 ;
   RECT 23.18 34.2 695.02 35.91 ;
   RECT 23.18 35.91 695.02 37.62 ;
   RECT 23.18 37.62 695.02 39.33 ;
   RECT 23.18 39.33 695.02 41.04 ;
   RECT 23.18 41.04 695.02 42.75 ;
   RECT 23.18 42.75 695.02 44.46 ;
   RECT 23.18 44.46 695.02 46.17 ;
   RECT 23.18 46.17 695.02 47.88 ;
   RECT 23.18 47.88 695.02 49.59 ;
   RECT 23.18 49.59 695.02 51.3 ;
   RECT 23.18 51.3 695.02 53.01 ;
   RECT 23.18 53.01 695.02 54.72 ;
   RECT 23.18 54.72 695.02 56.43 ;
   RECT 23.18 56.43 695.02 58.14 ;
   RECT 23.18 58.14 695.02 59.85 ;
   RECT 23.18 59.85 695.02 61.56 ;
   RECT 23.18 61.56 695.02 63.27 ;
   RECT 23.18 63.27 695.02 64.98 ;
   RECT 23.18 64.98 695.02 66.69 ;
   RECT 23.18 66.69 695.02 68.4 ;
   RECT 23.18 68.4 695.02 70.11 ;
   RECT 23.18 70.11 695.02 71.82 ;
   RECT 23.18 71.82 695.02 73.53 ;
   RECT 23.18 73.53 695.02 75.24 ;
   RECT 23.18 75.24 695.02 76.95 ;
   RECT 23.18 76.95 695.02 78.66 ;
   RECT 23.18 78.66 695.02 80.37 ;
   RECT 23.18 80.37 695.02 82.08 ;
   RECT 23.18 82.08 695.02 83.79 ;
   RECT 23.18 83.79 695.02 85.5 ;
   RECT 23.18 85.5 695.02 87.21 ;
   RECT 23.18 87.21 695.02 88.92 ;
   RECT 23.18 88.92 695.02 90.63 ;
   RECT 23.18 90.63 695.02 92.34 ;
   RECT 23.18 92.34 695.02 94.05 ;
   RECT 23.18 94.05 695.02 95.76 ;
   RECT 23.18 95.76 695.02 97.47 ;
   RECT 23.18 97.47 695.02 99.18 ;
   RECT 23.18 99.18 695.02 100.89 ;
   RECT 23.18 100.89 695.02 102.6 ;
   RECT 23.18 102.6 695.02 104.31 ;
   RECT 23.18 104.31 695.02 106.02 ;
   RECT 23.18 106.02 695.02 107.73 ;
   RECT 23.18 107.73 695.02 109.44 ;
   RECT 23.18 109.44 695.02 111.15 ;
   RECT 23.18 111.15 695.02 112.86 ;
   RECT 23.18 112.86 695.02 114.57 ;
   RECT 23.18 114.57 695.02 116.28 ;
   RECT 23.18 116.28 695.02 117.99 ;
   RECT 23.18 117.99 695.02 119.7 ;
   RECT 23.18 119.7 695.02 121.41 ;
   RECT 23.18 121.41 695.02 123.12 ;
   RECT 23.18 123.12 695.02 124.83 ;
   RECT 23.18 124.83 695.02 126.54 ;
   RECT 23.18 126.54 695.02 128.25 ;
   RECT 23.18 128.25 695.02 129.96 ;
   RECT 23.18 129.96 695.02 131.67 ;
   RECT 23.18 131.67 695.02 133.38 ;
   RECT 23.18 133.38 695.02 135.09 ;
   RECT 23.18 135.09 695.02 136.8 ;
   RECT 23.18 136.8 695.02 138.51 ;
   RECT 23.18 138.51 695.02 140.22 ;
   RECT 23.18 140.22 695.02 141.93 ;
   RECT 23.18 141.93 695.02 143.64 ;
   RECT 23.18 143.64 695.02 145.35 ;
   RECT 23.18 145.35 695.02 147.06 ;
   RECT 23.18 147.06 695.02 148.77 ;
   RECT 23.18 148.77 695.02 150.48 ;
   RECT 23.18 150.48 695.02 152.19 ;
   RECT 23.18 152.19 695.02 153.9 ;
   RECT 23.18 153.9 695.02 155.61 ;
   RECT 23.18 155.61 695.02 157.32 ;
   RECT 23.18 157.32 695.02 159.03 ;
   RECT 23.18 159.03 695.02 160.74 ;
   RECT 23.18 160.74 695.02 162.45 ;
   RECT 23.18 162.45 695.02 164.16 ;
   RECT 23.18 164.16 695.02 165.87 ;
   RECT 23.18 165.87 695.02 167.58 ;
   RECT 23.18 167.58 695.02 169.29 ;
   RECT 23.18 169.29 695.02 171.0 ;
   RECT 23.18 171.0 695.02 172.71 ;
   RECT 23.18 172.71 695.02 174.42 ;
   RECT 23.18 174.42 695.02 176.13 ;
   RECT 23.18 176.13 695.02 177.84 ;
   RECT 23.18 177.84 695.02 179.55 ;
   RECT 23.18 179.55 695.02 181.26 ;
   RECT 23.18 181.26 695.02 182.97 ;
   RECT 23.18 182.97 695.02 184.68 ;
   RECT 23.18 184.68 695.02 186.39 ;
   RECT 23.18 186.39 695.02 188.1 ;
   RECT 23.18 188.1 695.02 189.81 ;
   RECT 23.18 189.81 695.02 191.52 ;
   RECT 23.18 191.52 695.02 193.23 ;
   RECT 23.18 193.23 695.02 194.94 ;
   RECT 23.18 194.94 695.02 196.65 ;
   RECT 23.18 196.65 695.02 198.36 ;
   RECT 23.18 198.36 695.02 200.07 ;
   RECT 23.18 200.07 695.02 201.78 ;
   RECT 23.18 201.78 695.02 203.49 ;
   RECT 23.18 203.49 695.02 205.2 ;
   RECT 23.18 205.2 695.02 206.91 ;
   RECT 23.18 206.91 695.02 208.62 ;
   RECT 23.18 208.62 695.02 210.33 ;
   RECT 23.18 210.33 695.02 212.04 ;
   RECT 23.18 212.04 695.02 213.75 ;
   RECT 23.18 213.75 695.02 215.46 ;
   RECT 0.0 215.46 695.02 217.17 ;
   RECT 0.0 217.17 695.02 218.88 ;
   RECT 0.0 218.88 695.02 220.59 ;
   RECT 0.0 220.59 695.02 222.3 ;
   RECT 0.0 222.3 695.02 224.01 ;
   RECT 0.0 224.01 695.02 225.72 ;
   RECT 0.0 225.72 695.02 227.43 ;
   RECT 0.0 227.43 695.02 229.14 ;
   RECT 0.0 229.14 695.02 230.85 ;
   RECT 0.0 230.85 695.02 232.56 ;
   RECT 0.0 232.56 695.02 234.27 ;
   RECT 0.0 234.27 695.02 235.98 ;
   RECT 0.0 235.98 695.02 237.69 ;
   RECT 0.0 237.69 695.02 239.4 ;
   RECT 0.0 239.4 695.02 241.11 ;
   RECT 0.0 241.11 695.02 242.82 ;
   RECT 0.0 242.82 695.02 244.53 ;
   RECT 23.18 244.53 695.02 246.24 ;
   RECT 23.18 246.24 695.02 247.95 ;
   RECT 23.18 247.95 695.02 249.66 ;
   RECT 23.18 249.66 695.02 251.37 ;
   RECT 23.18 251.37 695.02 253.08 ;
   RECT 23.18 253.08 695.02 254.79 ;
   RECT 23.18 254.79 695.02 256.5 ;
   RECT 23.18 256.5 695.02 258.21 ;
   RECT 23.18 258.21 695.02 259.92 ;
   RECT 23.18 259.92 695.02 261.63 ;
   RECT 23.18 261.63 695.02 263.34 ;
   RECT 23.18 263.34 695.02 265.05 ;
   RECT 23.18 265.05 695.02 266.76 ;
   RECT 23.18 266.76 695.02 268.47 ;
   RECT 23.18 268.47 695.02 270.18 ;
   RECT 23.18 270.18 695.02 271.89 ;
   RECT 23.18 271.89 695.02 273.6 ;
   RECT 23.18 273.6 695.02 275.31 ;
   RECT 23.18 275.31 695.02 277.02 ;
   RECT 23.18 277.02 695.02 278.73 ;
   RECT 23.18 278.73 695.02 280.44 ;
   RECT 23.18 280.44 695.02 282.15 ;
   RECT 23.18 282.15 695.02 283.86 ;
   RECT 23.18 283.86 695.02 285.57 ;
   RECT 23.18 285.57 695.02 287.28 ;
   RECT 23.18 287.28 695.02 288.99 ;
   RECT 23.18 288.99 695.02 290.7 ;
   RECT 23.18 290.7 695.02 292.41 ;
   RECT 23.18 292.41 695.02 294.12 ;
   RECT 23.18 294.12 695.02 295.83 ;
   RECT 23.18 295.83 695.02 297.54 ;
   RECT 23.18 297.54 695.02 299.25 ;
   RECT 23.18 299.25 695.02 300.96 ;
   RECT 23.18 300.96 695.02 302.67 ;
   RECT 23.18 302.67 695.02 304.38 ;
   RECT 23.18 304.38 695.02 306.09 ;
   RECT 23.18 306.09 695.02 307.8 ;
   RECT 23.18 307.8 695.02 309.51 ;
   RECT 23.18 309.51 695.02 311.22 ;
   RECT 23.18 311.22 695.02 312.93 ;
   RECT 23.18 312.93 695.02 314.64 ;
   RECT 23.18 314.64 695.02 316.35 ;
   RECT 23.18 316.35 695.02 318.06 ;
   RECT 23.18 318.06 695.02 319.77 ;
   RECT 23.18 319.77 695.02 321.48 ;
   RECT 23.18 321.48 695.02 323.19 ;
   RECT 23.18 323.19 695.02 324.9 ;
   RECT 23.18 324.9 695.02 326.61 ;
   RECT 23.18 326.61 695.02 328.32 ;
   RECT 23.18 328.32 695.02 330.03 ;
   RECT 23.18 330.03 695.02 331.74 ;
   RECT 23.18 331.74 695.02 333.45 ;
   RECT 23.18 333.45 695.02 335.16 ;
   RECT 23.18 335.16 695.02 336.87 ;
   RECT 23.18 336.87 695.02 338.58 ;
   RECT 23.18 338.58 695.02 340.29 ;
   RECT 23.18 340.29 695.02 342.0 ;
   RECT 23.18 342.0 695.02 343.71 ;
   RECT 23.18 343.71 695.02 345.42 ;
   RECT 23.18 345.42 695.02 347.13 ;
   RECT 23.18 347.13 695.02 348.84 ;
   RECT 23.18 348.84 695.02 350.55 ;
   RECT 23.18 350.55 695.02 352.26 ;
   RECT 23.18 352.26 695.02 353.97 ;
   RECT 23.18 353.97 695.02 355.68 ;
   RECT 23.18 355.68 695.02 357.39 ;
   RECT 23.18 357.39 695.02 359.1 ;
   RECT 23.18 359.1 695.02 360.81 ;
   RECT 23.18 360.81 695.02 362.52 ;
   RECT 23.18 362.52 695.02 364.23 ;
   RECT 23.18 364.23 695.02 365.94 ;
   RECT 23.18 365.94 695.02 367.65 ;
   RECT 23.18 367.65 695.02 369.36 ;
   RECT 23.18 369.36 695.02 371.07 ;
   RECT 23.18 371.07 695.02 372.78 ;
   RECT 23.18 372.78 695.02 374.49 ;
   RECT 23.18 374.49 695.02 376.2 ;
   RECT 23.18 376.2 695.02 377.91 ;
   RECT 23.18 377.91 695.02 379.62 ;
   RECT 23.18 379.62 695.02 381.33 ;
   RECT 23.18 381.33 695.02 383.04 ;
   RECT 23.18 383.04 695.02 384.75 ;
   RECT 23.18 384.75 695.02 386.46 ;
   RECT 23.18 386.46 695.02 388.17 ;
   RECT 23.18 388.17 695.02 389.88 ;
   RECT 23.18 389.88 695.02 391.59 ;
   RECT 23.18 391.59 695.02 393.3 ;
   RECT 23.18 393.3 695.02 395.01 ;
   RECT 23.18 395.01 695.02 396.72 ;
   RECT 23.18 396.72 695.02 398.43 ;
   RECT 23.18 398.43 695.02 400.14 ;
   RECT 23.18 400.14 695.02 401.85 ;
   RECT 23.18 401.85 695.02 403.56 ;
   RECT 23.18 403.56 695.02 405.27 ;
   RECT 23.18 405.27 695.02 406.98 ;
   RECT 23.18 406.98 695.02 408.69 ;
   RECT 23.18 408.69 695.02 410.4 ;
   RECT 23.18 410.4 695.02 412.11 ;
   RECT 23.18 412.11 695.02 413.82 ;
   RECT 23.18 413.82 695.02 415.53 ;
   RECT 23.18 415.53 695.02 417.24 ;
   RECT 23.18 417.24 695.02 418.95 ;
   RECT 23.18 418.95 695.02 420.66 ;
   RECT 23.18 420.66 695.02 422.37 ;
   RECT 23.18 422.37 695.02 424.08 ;
   RECT 23.18 424.08 695.02 425.79 ;
   RECT 23.18 425.79 695.02 427.5 ;
   RECT 23.18 427.5 695.02 429.21 ;
   RECT 23.18 429.21 695.02 430.92 ;
   RECT 23.18 430.92 695.02 432.63 ;
   RECT 23.18 432.63 695.02 434.34 ;
   RECT 23.18 434.34 695.02 436.05 ;
   RECT 23.18 436.05 695.02 437.76 ;
   RECT 23.18 437.76 695.02 439.47 ;
   RECT 23.18 439.47 695.02 441.18 ;
   RECT 23.18 441.18 695.02 442.89 ;
   RECT 23.18 442.89 695.02 444.6 ;
   RECT 23.18 444.6 695.02 446.31 ;
   RECT 23.18 446.31 695.02 448.02 ;
   RECT 23.18 448.02 695.02 449.73 ;
   RECT 23.18 449.73 695.02 451.44 ;
   RECT 23.18 451.44 695.02 453.15 ;
   RECT 23.18 453.15 695.02 454.86 ;
   RECT 23.18 454.86 695.02 456.57 ;
   RECT 23.18 456.57 695.02 458.28 ;
   RECT 23.18 458.28 695.02 459.99 ;
   RECT 23.18 459.99 695.02 461.7 ;
   RECT 23.18 461.7 695.02 463.41 ;
   RECT 23.18 463.41 695.02 465.12 ;
   RECT 23.18 465.12 695.02 466.83 ;
   RECT 23.18 466.83 695.02 468.54 ;
   RECT 23.18 468.54 695.02 470.25 ;
   RECT 23.18 470.25 695.02 471.96 ;
   RECT 23.18 471.96 695.02 473.67 ;
   RECT 23.18 473.67 695.02 475.38 ;
  LAYER via3 ;
   RECT 23.18 0.0 695.02 1.71 ;
   RECT 23.18 1.71 695.02 3.42 ;
   RECT 23.18 3.42 695.02 5.13 ;
   RECT 23.18 5.13 695.02 6.84 ;
   RECT 23.18 6.84 695.02 8.55 ;
   RECT 23.18 8.55 695.02 10.26 ;
   RECT 23.18 10.26 695.02 11.97 ;
   RECT 23.18 11.97 695.02 13.68 ;
   RECT 23.18 13.68 695.02 15.39 ;
   RECT 23.18 15.39 695.02 17.1 ;
   RECT 23.18 17.1 695.02 18.81 ;
   RECT 23.18 18.81 695.02 20.52 ;
   RECT 23.18 20.52 695.02 22.23 ;
   RECT 23.18 22.23 695.02 23.94 ;
   RECT 23.18 23.94 695.02 25.65 ;
   RECT 23.18 25.65 695.02 27.36 ;
   RECT 23.18 27.36 695.02 29.07 ;
   RECT 23.18 29.07 695.02 30.78 ;
   RECT 23.18 30.78 695.02 32.49 ;
   RECT 23.18 32.49 695.02 34.2 ;
   RECT 23.18 34.2 695.02 35.91 ;
   RECT 23.18 35.91 695.02 37.62 ;
   RECT 23.18 37.62 695.02 39.33 ;
   RECT 23.18 39.33 695.02 41.04 ;
   RECT 23.18 41.04 695.02 42.75 ;
   RECT 23.18 42.75 695.02 44.46 ;
   RECT 23.18 44.46 695.02 46.17 ;
   RECT 23.18 46.17 695.02 47.88 ;
   RECT 23.18 47.88 695.02 49.59 ;
   RECT 23.18 49.59 695.02 51.3 ;
   RECT 23.18 51.3 695.02 53.01 ;
   RECT 23.18 53.01 695.02 54.72 ;
   RECT 23.18 54.72 695.02 56.43 ;
   RECT 23.18 56.43 695.02 58.14 ;
   RECT 23.18 58.14 695.02 59.85 ;
   RECT 23.18 59.85 695.02 61.56 ;
   RECT 23.18 61.56 695.02 63.27 ;
   RECT 23.18 63.27 695.02 64.98 ;
   RECT 23.18 64.98 695.02 66.69 ;
   RECT 23.18 66.69 695.02 68.4 ;
   RECT 23.18 68.4 695.02 70.11 ;
   RECT 23.18 70.11 695.02 71.82 ;
   RECT 23.18 71.82 695.02 73.53 ;
   RECT 23.18 73.53 695.02 75.24 ;
   RECT 23.18 75.24 695.02 76.95 ;
   RECT 23.18 76.95 695.02 78.66 ;
   RECT 23.18 78.66 695.02 80.37 ;
   RECT 23.18 80.37 695.02 82.08 ;
   RECT 23.18 82.08 695.02 83.79 ;
   RECT 23.18 83.79 695.02 85.5 ;
   RECT 23.18 85.5 695.02 87.21 ;
   RECT 23.18 87.21 695.02 88.92 ;
   RECT 23.18 88.92 695.02 90.63 ;
   RECT 23.18 90.63 695.02 92.34 ;
   RECT 23.18 92.34 695.02 94.05 ;
   RECT 23.18 94.05 695.02 95.76 ;
   RECT 23.18 95.76 695.02 97.47 ;
   RECT 23.18 97.47 695.02 99.18 ;
   RECT 23.18 99.18 695.02 100.89 ;
   RECT 23.18 100.89 695.02 102.6 ;
   RECT 23.18 102.6 695.02 104.31 ;
   RECT 23.18 104.31 695.02 106.02 ;
   RECT 23.18 106.02 695.02 107.73 ;
   RECT 23.18 107.73 695.02 109.44 ;
   RECT 23.18 109.44 695.02 111.15 ;
   RECT 23.18 111.15 695.02 112.86 ;
   RECT 23.18 112.86 695.02 114.57 ;
   RECT 23.18 114.57 695.02 116.28 ;
   RECT 23.18 116.28 695.02 117.99 ;
   RECT 23.18 117.99 695.02 119.7 ;
   RECT 23.18 119.7 695.02 121.41 ;
   RECT 23.18 121.41 695.02 123.12 ;
   RECT 23.18 123.12 695.02 124.83 ;
   RECT 23.18 124.83 695.02 126.54 ;
   RECT 23.18 126.54 695.02 128.25 ;
   RECT 23.18 128.25 695.02 129.96 ;
   RECT 23.18 129.96 695.02 131.67 ;
   RECT 23.18 131.67 695.02 133.38 ;
   RECT 23.18 133.38 695.02 135.09 ;
   RECT 23.18 135.09 695.02 136.8 ;
   RECT 23.18 136.8 695.02 138.51 ;
   RECT 23.18 138.51 695.02 140.22 ;
   RECT 23.18 140.22 695.02 141.93 ;
   RECT 23.18 141.93 695.02 143.64 ;
   RECT 23.18 143.64 695.02 145.35 ;
   RECT 23.18 145.35 695.02 147.06 ;
   RECT 23.18 147.06 695.02 148.77 ;
   RECT 23.18 148.77 695.02 150.48 ;
   RECT 23.18 150.48 695.02 152.19 ;
   RECT 23.18 152.19 695.02 153.9 ;
   RECT 23.18 153.9 695.02 155.61 ;
   RECT 23.18 155.61 695.02 157.32 ;
   RECT 23.18 157.32 695.02 159.03 ;
   RECT 23.18 159.03 695.02 160.74 ;
   RECT 23.18 160.74 695.02 162.45 ;
   RECT 23.18 162.45 695.02 164.16 ;
   RECT 23.18 164.16 695.02 165.87 ;
   RECT 23.18 165.87 695.02 167.58 ;
   RECT 23.18 167.58 695.02 169.29 ;
   RECT 23.18 169.29 695.02 171.0 ;
   RECT 23.18 171.0 695.02 172.71 ;
   RECT 23.18 172.71 695.02 174.42 ;
   RECT 23.18 174.42 695.02 176.13 ;
   RECT 23.18 176.13 695.02 177.84 ;
   RECT 23.18 177.84 695.02 179.55 ;
   RECT 23.18 179.55 695.02 181.26 ;
   RECT 23.18 181.26 695.02 182.97 ;
   RECT 23.18 182.97 695.02 184.68 ;
   RECT 23.18 184.68 695.02 186.39 ;
   RECT 23.18 186.39 695.02 188.1 ;
   RECT 23.18 188.1 695.02 189.81 ;
   RECT 23.18 189.81 695.02 191.52 ;
   RECT 23.18 191.52 695.02 193.23 ;
   RECT 23.18 193.23 695.02 194.94 ;
   RECT 23.18 194.94 695.02 196.65 ;
   RECT 23.18 196.65 695.02 198.36 ;
   RECT 23.18 198.36 695.02 200.07 ;
   RECT 23.18 200.07 695.02 201.78 ;
   RECT 23.18 201.78 695.02 203.49 ;
   RECT 23.18 203.49 695.02 205.2 ;
   RECT 23.18 205.2 695.02 206.91 ;
   RECT 23.18 206.91 695.02 208.62 ;
   RECT 23.18 208.62 695.02 210.33 ;
   RECT 23.18 210.33 695.02 212.04 ;
   RECT 23.18 212.04 695.02 213.75 ;
   RECT 23.18 213.75 695.02 215.46 ;
   RECT 0.0 215.46 695.02 217.17 ;
   RECT 0.0 217.17 695.02 218.88 ;
   RECT 0.0 218.88 695.02 220.59 ;
   RECT 0.0 220.59 695.02 222.3 ;
   RECT 0.0 222.3 695.02 224.01 ;
   RECT 0.0 224.01 695.02 225.72 ;
   RECT 0.0 225.72 695.02 227.43 ;
   RECT 0.0 227.43 695.02 229.14 ;
   RECT 0.0 229.14 695.02 230.85 ;
   RECT 0.0 230.85 695.02 232.56 ;
   RECT 0.0 232.56 695.02 234.27 ;
   RECT 0.0 234.27 695.02 235.98 ;
   RECT 0.0 235.98 695.02 237.69 ;
   RECT 0.0 237.69 695.02 239.4 ;
   RECT 0.0 239.4 695.02 241.11 ;
   RECT 0.0 241.11 695.02 242.82 ;
   RECT 0.0 242.82 695.02 244.53 ;
   RECT 23.18 244.53 695.02 246.24 ;
   RECT 23.18 246.24 695.02 247.95 ;
   RECT 23.18 247.95 695.02 249.66 ;
   RECT 23.18 249.66 695.02 251.37 ;
   RECT 23.18 251.37 695.02 253.08 ;
   RECT 23.18 253.08 695.02 254.79 ;
   RECT 23.18 254.79 695.02 256.5 ;
   RECT 23.18 256.5 695.02 258.21 ;
   RECT 23.18 258.21 695.02 259.92 ;
   RECT 23.18 259.92 695.02 261.63 ;
   RECT 23.18 261.63 695.02 263.34 ;
   RECT 23.18 263.34 695.02 265.05 ;
   RECT 23.18 265.05 695.02 266.76 ;
   RECT 23.18 266.76 695.02 268.47 ;
   RECT 23.18 268.47 695.02 270.18 ;
   RECT 23.18 270.18 695.02 271.89 ;
   RECT 23.18 271.89 695.02 273.6 ;
   RECT 23.18 273.6 695.02 275.31 ;
   RECT 23.18 275.31 695.02 277.02 ;
   RECT 23.18 277.02 695.02 278.73 ;
   RECT 23.18 278.73 695.02 280.44 ;
   RECT 23.18 280.44 695.02 282.15 ;
   RECT 23.18 282.15 695.02 283.86 ;
   RECT 23.18 283.86 695.02 285.57 ;
   RECT 23.18 285.57 695.02 287.28 ;
   RECT 23.18 287.28 695.02 288.99 ;
   RECT 23.18 288.99 695.02 290.7 ;
   RECT 23.18 290.7 695.02 292.41 ;
   RECT 23.18 292.41 695.02 294.12 ;
   RECT 23.18 294.12 695.02 295.83 ;
   RECT 23.18 295.83 695.02 297.54 ;
   RECT 23.18 297.54 695.02 299.25 ;
   RECT 23.18 299.25 695.02 300.96 ;
   RECT 23.18 300.96 695.02 302.67 ;
   RECT 23.18 302.67 695.02 304.38 ;
   RECT 23.18 304.38 695.02 306.09 ;
   RECT 23.18 306.09 695.02 307.8 ;
   RECT 23.18 307.8 695.02 309.51 ;
   RECT 23.18 309.51 695.02 311.22 ;
   RECT 23.18 311.22 695.02 312.93 ;
   RECT 23.18 312.93 695.02 314.64 ;
   RECT 23.18 314.64 695.02 316.35 ;
   RECT 23.18 316.35 695.02 318.06 ;
   RECT 23.18 318.06 695.02 319.77 ;
   RECT 23.18 319.77 695.02 321.48 ;
   RECT 23.18 321.48 695.02 323.19 ;
   RECT 23.18 323.19 695.02 324.9 ;
   RECT 23.18 324.9 695.02 326.61 ;
   RECT 23.18 326.61 695.02 328.32 ;
   RECT 23.18 328.32 695.02 330.03 ;
   RECT 23.18 330.03 695.02 331.74 ;
   RECT 23.18 331.74 695.02 333.45 ;
   RECT 23.18 333.45 695.02 335.16 ;
   RECT 23.18 335.16 695.02 336.87 ;
   RECT 23.18 336.87 695.02 338.58 ;
   RECT 23.18 338.58 695.02 340.29 ;
   RECT 23.18 340.29 695.02 342.0 ;
   RECT 23.18 342.0 695.02 343.71 ;
   RECT 23.18 343.71 695.02 345.42 ;
   RECT 23.18 345.42 695.02 347.13 ;
   RECT 23.18 347.13 695.02 348.84 ;
   RECT 23.18 348.84 695.02 350.55 ;
   RECT 23.18 350.55 695.02 352.26 ;
   RECT 23.18 352.26 695.02 353.97 ;
   RECT 23.18 353.97 695.02 355.68 ;
   RECT 23.18 355.68 695.02 357.39 ;
   RECT 23.18 357.39 695.02 359.1 ;
   RECT 23.18 359.1 695.02 360.81 ;
   RECT 23.18 360.81 695.02 362.52 ;
   RECT 23.18 362.52 695.02 364.23 ;
   RECT 23.18 364.23 695.02 365.94 ;
   RECT 23.18 365.94 695.02 367.65 ;
   RECT 23.18 367.65 695.02 369.36 ;
   RECT 23.18 369.36 695.02 371.07 ;
   RECT 23.18 371.07 695.02 372.78 ;
   RECT 23.18 372.78 695.02 374.49 ;
   RECT 23.18 374.49 695.02 376.2 ;
   RECT 23.18 376.2 695.02 377.91 ;
   RECT 23.18 377.91 695.02 379.62 ;
   RECT 23.18 379.62 695.02 381.33 ;
   RECT 23.18 381.33 695.02 383.04 ;
   RECT 23.18 383.04 695.02 384.75 ;
   RECT 23.18 384.75 695.02 386.46 ;
   RECT 23.18 386.46 695.02 388.17 ;
   RECT 23.18 388.17 695.02 389.88 ;
   RECT 23.18 389.88 695.02 391.59 ;
   RECT 23.18 391.59 695.02 393.3 ;
   RECT 23.18 393.3 695.02 395.01 ;
   RECT 23.18 395.01 695.02 396.72 ;
   RECT 23.18 396.72 695.02 398.43 ;
   RECT 23.18 398.43 695.02 400.14 ;
   RECT 23.18 400.14 695.02 401.85 ;
   RECT 23.18 401.85 695.02 403.56 ;
   RECT 23.18 403.56 695.02 405.27 ;
   RECT 23.18 405.27 695.02 406.98 ;
   RECT 23.18 406.98 695.02 408.69 ;
   RECT 23.18 408.69 695.02 410.4 ;
   RECT 23.18 410.4 695.02 412.11 ;
   RECT 23.18 412.11 695.02 413.82 ;
   RECT 23.18 413.82 695.02 415.53 ;
   RECT 23.18 415.53 695.02 417.24 ;
   RECT 23.18 417.24 695.02 418.95 ;
   RECT 23.18 418.95 695.02 420.66 ;
   RECT 23.18 420.66 695.02 422.37 ;
   RECT 23.18 422.37 695.02 424.08 ;
   RECT 23.18 424.08 695.02 425.79 ;
   RECT 23.18 425.79 695.02 427.5 ;
   RECT 23.18 427.5 695.02 429.21 ;
   RECT 23.18 429.21 695.02 430.92 ;
   RECT 23.18 430.92 695.02 432.63 ;
   RECT 23.18 432.63 695.02 434.34 ;
   RECT 23.18 434.34 695.02 436.05 ;
   RECT 23.18 436.05 695.02 437.76 ;
   RECT 23.18 437.76 695.02 439.47 ;
   RECT 23.18 439.47 695.02 441.18 ;
   RECT 23.18 441.18 695.02 442.89 ;
   RECT 23.18 442.89 695.02 444.6 ;
   RECT 23.18 444.6 695.02 446.31 ;
   RECT 23.18 446.31 695.02 448.02 ;
   RECT 23.18 448.02 695.02 449.73 ;
   RECT 23.18 449.73 695.02 451.44 ;
   RECT 23.18 451.44 695.02 453.15 ;
   RECT 23.18 453.15 695.02 454.86 ;
   RECT 23.18 454.86 695.02 456.57 ;
   RECT 23.18 456.57 695.02 458.28 ;
   RECT 23.18 458.28 695.02 459.99 ;
   RECT 23.18 459.99 695.02 461.7 ;
   RECT 23.18 461.7 695.02 463.41 ;
   RECT 23.18 463.41 695.02 465.12 ;
   RECT 23.18 465.12 695.02 466.83 ;
   RECT 23.18 466.83 695.02 468.54 ;
   RECT 23.18 468.54 695.02 470.25 ;
   RECT 23.18 470.25 695.02 471.96 ;
   RECT 23.18 471.96 695.02 473.67 ;
   RECT 23.18 473.67 695.02 475.38 ;
  LAYER metal4 ;
   RECT 23.18 0.0 695.02 1.71 ;
   RECT 23.18 1.71 695.02 3.42 ;
   RECT 23.18 3.42 695.02 5.13 ;
   RECT 23.18 5.13 695.02 6.84 ;
   RECT 23.18 6.84 695.02 8.55 ;
   RECT 23.18 8.55 695.02 10.26 ;
   RECT 23.18 10.26 695.02 11.97 ;
   RECT 23.18 11.97 695.02 13.68 ;
   RECT 23.18 13.68 695.02 15.39 ;
   RECT 23.18 15.39 695.02 17.1 ;
   RECT 23.18 17.1 695.02 18.81 ;
   RECT 23.18 18.81 695.02 20.52 ;
   RECT 23.18 20.52 695.02 22.23 ;
   RECT 23.18 22.23 695.02 23.94 ;
   RECT 23.18 23.94 695.02 25.65 ;
   RECT 23.18 25.65 695.02 27.36 ;
   RECT 23.18 27.36 695.02 29.07 ;
   RECT 23.18 29.07 695.02 30.78 ;
   RECT 23.18 30.78 695.02 32.49 ;
   RECT 23.18 32.49 695.02 34.2 ;
   RECT 23.18 34.2 695.02 35.91 ;
   RECT 23.18 35.91 695.02 37.62 ;
   RECT 23.18 37.62 695.02 39.33 ;
   RECT 23.18 39.33 695.02 41.04 ;
   RECT 23.18 41.04 695.02 42.75 ;
   RECT 23.18 42.75 695.02 44.46 ;
   RECT 23.18 44.46 695.02 46.17 ;
   RECT 23.18 46.17 695.02 47.88 ;
   RECT 23.18 47.88 695.02 49.59 ;
   RECT 23.18 49.59 695.02 51.3 ;
   RECT 23.18 51.3 695.02 53.01 ;
   RECT 23.18 53.01 695.02 54.72 ;
   RECT 23.18 54.72 695.02 56.43 ;
   RECT 23.18 56.43 695.02 58.14 ;
   RECT 23.18 58.14 695.02 59.85 ;
   RECT 23.18 59.85 695.02 61.56 ;
   RECT 23.18 61.56 695.02 63.27 ;
   RECT 23.18 63.27 695.02 64.98 ;
   RECT 23.18 64.98 695.02 66.69 ;
   RECT 23.18 66.69 695.02 68.4 ;
   RECT 23.18 68.4 695.02 70.11 ;
   RECT 23.18 70.11 695.02 71.82 ;
   RECT 23.18 71.82 695.02 73.53 ;
   RECT 23.18 73.53 695.02 75.24 ;
   RECT 23.18 75.24 695.02 76.95 ;
   RECT 23.18 76.95 695.02 78.66 ;
   RECT 23.18 78.66 695.02 80.37 ;
   RECT 23.18 80.37 695.02 82.08 ;
   RECT 23.18 82.08 695.02 83.79 ;
   RECT 23.18 83.79 695.02 85.5 ;
   RECT 23.18 85.5 695.02 87.21 ;
   RECT 23.18 87.21 695.02 88.92 ;
   RECT 23.18 88.92 695.02 90.63 ;
   RECT 23.18 90.63 695.02 92.34 ;
   RECT 23.18 92.34 695.02 94.05 ;
   RECT 23.18 94.05 695.02 95.76 ;
   RECT 23.18 95.76 695.02 97.47 ;
   RECT 23.18 97.47 695.02 99.18 ;
   RECT 23.18 99.18 695.02 100.89 ;
   RECT 23.18 100.89 695.02 102.6 ;
   RECT 23.18 102.6 695.02 104.31 ;
   RECT 23.18 104.31 695.02 106.02 ;
   RECT 23.18 106.02 695.02 107.73 ;
   RECT 23.18 107.73 695.02 109.44 ;
   RECT 23.18 109.44 695.02 111.15 ;
   RECT 23.18 111.15 695.02 112.86 ;
   RECT 23.18 112.86 695.02 114.57 ;
   RECT 23.18 114.57 695.02 116.28 ;
   RECT 23.18 116.28 695.02 117.99 ;
   RECT 23.18 117.99 695.02 119.7 ;
   RECT 23.18 119.7 695.02 121.41 ;
   RECT 23.18 121.41 695.02 123.12 ;
   RECT 23.18 123.12 695.02 124.83 ;
   RECT 23.18 124.83 695.02 126.54 ;
   RECT 23.18 126.54 695.02 128.25 ;
   RECT 23.18 128.25 695.02 129.96 ;
   RECT 23.18 129.96 695.02 131.67 ;
   RECT 23.18 131.67 695.02 133.38 ;
   RECT 23.18 133.38 695.02 135.09 ;
   RECT 23.18 135.09 695.02 136.8 ;
   RECT 23.18 136.8 695.02 138.51 ;
   RECT 23.18 138.51 695.02 140.22 ;
   RECT 23.18 140.22 695.02 141.93 ;
   RECT 23.18 141.93 695.02 143.64 ;
   RECT 23.18 143.64 695.02 145.35 ;
   RECT 23.18 145.35 695.02 147.06 ;
   RECT 23.18 147.06 695.02 148.77 ;
   RECT 23.18 148.77 695.02 150.48 ;
   RECT 23.18 150.48 695.02 152.19 ;
   RECT 23.18 152.19 695.02 153.9 ;
   RECT 23.18 153.9 695.02 155.61 ;
   RECT 23.18 155.61 695.02 157.32 ;
   RECT 23.18 157.32 695.02 159.03 ;
   RECT 23.18 159.03 695.02 160.74 ;
   RECT 23.18 160.74 695.02 162.45 ;
   RECT 23.18 162.45 695.02 164.16 ;
   RECT 23.18 164.16 695.02 165.87 ;
   RECT 23.18 165.87 695.02 167.58 ;
   RECT 23.18 167.58 695.02 169.29 ;
   RECT 23.18 169.29 695.02 171.0 ;
   RECT 23.18 171.0 695.02 172.71 ;
   RECT 23.18 172.71 695.02 174.42 ;
   RECT 23.18 174.42 695.02 176.13 ;
   RECT 23.18 176.13 695.02 177.84 ;
   RECT 23.18 177.84 695.02 179.55 ;
   RECT 23.18 179.55 695.02 181.26 ;
   RECT 23.18 181.26 695.02 182.97 ;
   RECT 23.18 182.97 695.02 184.68 ;
   RECT 23.18 184.68 695.02 186.39 ;
   RECT 23.18 186.39 695.02 188.1 ;
   RECT 23.18 188.1 695.02 189.81 ;
   RECT 23.18 189.81 695.02 191.52 ;
   RECT 23.18 191.52 695.02 193.23 ;
   RECT 23.18 193.23 695.02 194.94 ;
   RECT 23.18 194.94 695.02 196.65 ;
   RECT 23.18 196.65 695.02 198.36 ;
   RECT 23.18 198.36 695.02 200.07 ;
   RECT 23.18 200.07 695.02 201.78 ;
   RECT 23.18 201.78 695.02 203.49 ;
   RECT 23.18 203.49 695.02 205.2 ;
   RECT 23.18 205.2 695.02 206.91 ;
   RECT 23.18 206.91 695.02 208.62 ;
   RECT 23.18 208.62 695.02 210.33 ;
   RECT 23.18 210.33 695.02 212.04 ;
   RECT 23.18 212.04 695.02 213.75 ;
   RECT 23.18 213.75 695.02 215.46 ;
   RECT 0.0 215.46 695.02 217.17 ;
   RECT 0.0 217.17 695.02 218.88 ;
   RECT 0.0 218.88 695.02 220.59 ;
   RECT 0.0 220.59 695.02 222.3 ;
   RECT 0.0 222.3 695.02 224.01 ;
   RECT 0.0 224.01 695.02 225.72 ;
   RECT 0.0 225.72 695.02 227.43 ;
   RECT 0.0 227.43 695.02 229.14 ;
   RECT 0.0 229.14 695.02 230.85 ;
   RECT 0.0 230.85 695.02 232.56 ;
   RECT 0.0 232.56 695.02 234.27 ;
   RECT 0.0 234.27 695.02 235.98 ;
   RECT 0.0 235.98 695.02 237.69 ;
   RECT 0.0 237.69 695.02 239.4 ;
   RECT 0.0 239.4 695.02 241.11 ;
   RECT 0.0 241.11 695.02 242.82 ;
   RECT 0.0 242.82 695.02 244.53 ;
   RECT 23.18 244.53 695.02 246.24 ;
   RECT 23.18 246.24 695.02 247.95 ;
   RECT 23.18 247.95 695.02 249.66 ;
   RECT 23.18 249.66 695.02 251.37 ;
   RECT 23.18 251.37 695.02 253.08 ;
   RECT 23.18 253.08 695.02 254.79 ;
   RECT 23.18 254.79 695.02 256.5 ;
   RECT 23.18 256.5 695.02 258.21 ;
   RECT 23.18 258.21 695.02 259.92 ;
   RECT 23.18 259.92 695.02 261.63 ;
   RECT 23.18 261.63 695.02 263.34 ;
   RECT 23.18 263.34 695.02 265.05 ;
   RECT 23.18 265.05 695.02 266.76 ;
   RECT 23.18 266.76 695.02 268.47 ;
   RECT 23.18 268.47 695.02 270.18 ;
   RECT 23.18 270.18 695.02 271.89 ;
   RECT 23.18 271.89 695.02 273.6 ;
   RECT 23.18 273.6 695.02 275.31 ;
   RECT 23.18 275.31 695.02 277.02 ;
   RECT 23.18 277.02 695.02 278.73 ;
   RECT 23.18 278.73 695.02 280.44 ;
   RECT 23.18 280.44 695.02 282.15 ;
   RECT 23.18 282.15 695.02 283.86 ;
   RECT 23.18 283.86 695.02 285.57 ;
   RECT 23.18 285.57 695.02 287.28 ;
   RECT 23.18 287.28 695.02 288.99 ;
   RECT 23.18 288.99 695.02 290.7 ;
   RECT 23.18 290.7 695.02 292.41 ;
   RECT 23.18 292.41 695.02 294.12 ;
   RECT 23.18 294.12 695.02 295.83 ;
   RECT 23.18 295.83 695.02 297.54 ;
   RECT 23.18 297.54 695.02 299.25 ;
   RECT 23.18 299.25 695.02 300.96 ;
   RECT 23.18 300.96 695.02 302.67 ;
   RECT 23.18 302.67 695.02 304.38 ;
   RECT 23.18 304.38 695.02 306.09 ;
   RECT 23.18 306.09 695.02 307.8 ;
   RECT 23.18 307.8 695.02 309.51 ;
   RECT 23.18 309.51 695.02 311.22 ;
   RECT 23.18 311.22 695.02 312.93 ;
   RECT 23.18 312.93 695.02 314.64 ;
   RECT 23.18 314.64 695.02 316.35 ;
   RECT 23.18 316.35 695.02 318.06 ;
   RECT 23.18 318.06 695.02 319.77 ;
   RECT 23.18 319.77 695.02 321.48 ;
   RECT 23.18 321.48 695.02 323.19 ;
   RECT 23.18 323.19 695.02 324.9 ;
   RECT 23.18 324.9 695.02 326.61 ;
   RECT 23.18 326.61 695.02 328.32 ;
   RECT 23.18 328.32 695.02 330.03 ;
   RECT 23.18 330.03 695.02 331.74 ;
   RECT 23.18 331.74 695.02 333.45 ;
   RECT 23.18 333.45 695.02 335.16 ;
   RECT 23.18 335.16 695.02 336.87 ;
   RECT 23.18 336.87 695.02 338.58 ;
   RECT 23.18 338.58 695.02 340.29 ;
   RECT 23.18 340.29 695.02 342.0 ;
   RECT 23.18 342.0 695.02 343.71 ;
   RECT 23.18 343.71 695.02 345.42 ;
   RECT 23.18 345.42 695.02 347.13 ;
   RECT 23.18 347.13 695.02 348.84 ;
   RECT 23.18 348.84 695.02 350.55 ;
   RECT 23.18 350.55 695.02 352.26 ;
   RECT 23.18 352.26 695.02 353.97 ;
   RECT 23.18 353.97 695.02 355.68 ;
   RECT 23.18 355.68 695.02 357.39 ;
   RECT 23.18 357.39 695.02 359.1 ;
   RECT 23.18 359.1 695.02 360.81 ;
   RECT 23.18 360.81 695.02 362.52 ;
   RECT 23.18 362.52 695.02 364.23 ;
   RECT 23.18 364.23 695.02 365.94 ;
   RECT 23.18 365.94 695.02 367.65 ;
   RECT 23.18 367.65 695.02 369.36 ;
   RECT 23.18 369.36 695.02 371.07 ;
   RECT 23.18 371.07 695.02 372.78 ;
   RECT 23.18 372.78 695.02 374.49 ;
   RECT 23.18 374.49 695.02 376.2 ;
   RECT 23.18 376.2 695.02 377.91 ;
   RECT 23.18 377.91 695.02 379.62 ;
   RECT 23.18 379.62 695.02 381.33 ;
   RECT 23.18 381.33 695.02 383.04 ;
   RECT 23.18 383.04 695.02 384.75 ;
   RECT 23.18 384.75 695.02 386.46 ;
   RECT 23.18 386.46 695.02 388.17 ;
   RECT 23.18 388.17 695.02 389.88 ;
   RECT 23.18 389.88 695.02 391.59 ;
   RECT 23.18 391.59 695.02 393.3 ;
   RECT 23.18 393.3 695.02 395.01 ;
   RECT 23.18 395.01 695.02 396.72 ;
   RECT 23.18 396.72 695.02 398.43 ;
   RECT 23.18 398.43 695.02 400.14 ;
   RECT 23.18 400.14 695.02 401.85 ;
   RECT 23.18 401.85 695.02 403.56 ;
   RECT 23.18 403.56 695.02 405.27 ;
   RECT 23.18 405.27 695.02 406.98 ;
   RECT 23.18 406.98 695.02 408.69 ;
   RECT 23.18 408.69 695.02 410.4 ;
   RECT 23.18 410.4 695.02 412.11 ;
   RECT 23.18 412.11 695.02 413.82 ;
   RECT 23.18 413.82 695.02 415.53 ;
   RECT 23.18 415.53 695.02 417.24 ;
   RECT 23.18 417.24 695.02 418.95 ;
   RECT 23.18 418.95 695.02 420.66 ;
   RECT 23.18 420.66 695.02 422.37 ;
   RECT 23.18 422.37 695.02 424.08 ;
   RECT 23.18 424.08 695.02 425.79 ;
   RECT 23.18 425.79 695.02 427.5 ;
   RECT 23.18 427.5 695.02 429.21 ;
   RECT 23.18 429.21 695.02 430.92 ;
   RECT 23.18 430.92 695.02 432.63 ;
   RECT 23.18 432.63 695.02 434.34 ;
   RECT 23.18 434.34 695.02 436.05 ;
   RECT 23.18 436.05 695.02 437.76 ;
   RECT 23.18 437.76 695.02 439.47 ;
   RECT 23.18 439.47 695.02 441.18 ;
   RECT 23.18 441.18 695.02 442.89 ;
   RECT 23.18 442.89 695.02 444.6 ;
   RECT 23.18 444.6 695.02 446.31 ;
   RECT 23.18 446.31 695.02 448.02 ;
   RECT 23.18 448.02 695.02 449.73 ;
   RECT 23.18 449.73 695.02 451.44 ;
   RECT 23.18 451.44 695.02 453.15 ;
   RECT 23.18 453.15 695.02 454.86 ;
   RECT 23.18 454.86 695.02 456.57 ;
   RECT 23.18 456.57 695.02 458.28 ;
   RECT 23.18 458.28 695.02 459.99 ;
   RECT 23.18 459.99 695.02 461.7 ;
   RECT 23.18 461.7 695.02 463.41 ;
   RECT 23.18 463.41 695.02 465.12 ;
   RECT 23.18 465.12 695.02 466.83 ;
   RECT 23.18 466.83 695.02 468.54 ;
   RECT 23.18 468.54 695.02 470.25 ;
   RECT 23.18 470.25 695.02 471.96 ;
   RECT 23.18 471.96 695.02 473.67 ;
   RECT 23.18 473.67 695.02 475.38 ;
 END
END block_1829x2502_263

MACRO block_1338x1773_192
 CLASS BLOCK ;
 FOREIGN block_1338x1773_192 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 508.44 BY 336.87 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 330.695 26.885 331.265 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 322.525 26.885 323.095 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 230.755 26.885 231.325 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 222.585 26.885 223.155 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 214.415 26.885 214.985 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 206.245 26.885 206.815 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 198.075 26.885 198.645 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 189.905 26.885 190.475 ;
  END
 END o7
 PIN o8
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 181.735 26.885 182.305 ;
  END
 END o8
 PIN o9
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 145.255 26.885 145.825 ;
  END
 END o9
 PIN o10
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 137.085 26.885 137.655 ;
  END
 END o10
 PIN o11
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 128.915 26.885 129.485 ;
  END
 END o11
 PIN o12
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 314.355 26.885 314.925 ;
  END
 END o12
 PIN o13
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 120.745 26.885 121.315 ;
  END
 END o13
 PIN o14
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 112.575 26.885 113.145 ;
  END
 END o14
 PIN o15
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 104.405 26.885 104.975 ;
  END
 END o15
 PIN o16
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 96.235 26.885 96.805 ;
  END
 END o16
 PIN o17
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 88.065 26.885 88.635 ;
  END
 END o17
 PIN o18
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 61.655 26.885 62.225 ;
  END
 END o18
 PIN o19
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 53.485 26.885 54.055 ;
  END
 END o19
 PIN o20
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 45.315 26.885 45.885 ;
  END
 END o20
 PIN o21
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 37.145 26.885 37.715 ;
  END
 END o21
 PIN o22
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 28.975 26.885 29.545 ;
  END
 END o22
 PIN o23
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 306.185 26.885 306.755 ;
  END
 END o23
 PIN o24
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 20.805 26.885 21.375 ;
  END
 END o24
 PIN o25
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 12.635 26.885 13.205 ;
  END
 END o25
 PIN o26
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 4.465 26.885 5.035 ;
  END
 END o26
 PIN o27
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 298.015 26.885 298.585 ;
  END
 END o27
 PIN o28
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 289.845 26.885 290.415 ;
  END
 END o28
 PIN o29
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 281.675 26.885 282.245 ;
  END
 END o29
 PIN o30
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 273.505 26.885 274.075 ;
  END
 END o30
 PIN o31
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 265.335 26.885 265.905 ;
  END
 END o31
 PIN o32
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 238.925 26.885 239.495 ;
  END
 END o32
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 174.705 3.705 175.275 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 153.045 3.705 153.615 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 157.605 3.705 158.175 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 169.385 3.705 169.955 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 165.015 3.705 165.585 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 174.325 4.465 174.895 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 175.085 4.465 175.655 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 175.465 3.705 176.035 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 165.775 3.705 166.345 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 152.665 4.465 153.235 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 157.985 4.465 158.555 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 161.215 3.705 161.785 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 158.365 3.705 158.935 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 156.275 3.705 156.845 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 153.805 3.705 154.375 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 152.285 3.705 152.855 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 13.015 175.845 13.585 176.415 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 14.155 175.845 14.725 176.415 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 13.015 162.545 13.585 163.115 ;
  END
 END i18
 PIN i19
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 14.155 162.545 14.725 163.115 ;
  END
 END i19
 PIN i20
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 332.405 26.885 332.975 ;
  END
 END i20
 PIN i21
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 324.235 26.885 324.805 ;
  END
 END i21
 PIN i22
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 232.465 26.885 233.035 ;
  END
 END i22
 PIN i23
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 224.295 26.885 224.865 ;
  END
 END i23
 PIN i24
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 216.125 26.885 216.695 ;
  END
 END i24
 PIN i25
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 207.955 26.885 208.525 ;
  END
 END i25
 PIN i26
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 199.785 26.885 200.355 ;
  END
 END i26
 PIN i27
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 191.615 26.885 192.185 ;
  END
 END i27
 PIN i28
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 183.445 26.885 184.015 ;
  END
 END i28
 PIN i29
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 143.545 26.885 144.115 ;
  END
 END i29
 PIN i30
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 135.375 26.885 135.945 ;
  END
 END i30
 PIN i31
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 127.205 26.885 127.775 ;
  END
 END i31
 PIN i32
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 316.065 26.885 316.635 ;
  END
 END i32
 PIN i33
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 119.035 26.885 119.605 ;
  END
 END i33
 PIN i34
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 110.865 26.885 111.435 ;
  END
 END i34
 PIN i35
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 102.695 26.885 103.265 ;
  END
 END i35
 PIN i36
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 94.525 26.885 95.095 ;
  END
 END i36
 PIN i37
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 86.355 26.885 86.925 ;
  END
 END i37
 PIN i38
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 59.945 26.885 60.515 ;
  END
 END i38
 PIN i39
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 51.775 26.885 52.345 ;
  END
 END i39
 PIN i40
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 43.605 26.885 44.175 ;
  END
 END i40
 PIN i41
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 35.435 26.885 36.005 ;
  END
 END i41
 PIN i42
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 27.265 26.885 27.835 ;
  END
 END i42
 PIN i43
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 307.895 26.885 308.465 ;
  END
 END i43
 PIN i44
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 19.095 26.885 19.665 ;
  END
 END i44
 PIN i45
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 10.925 26.885 11.495 ;
  END
 END i45
 PIN i46
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 2.755 26.885 3.325 ;
  END
 END i46
 PIN i47
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 299.725 26.885 300.295 ;
  END
 END i47
 PIN i48
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 291.555 26.885 292.125 ;
  END
 END i48
 PIN i49
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 283.385 26.885 283.955 ;
  END
 END i49
 PIN i50
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 275.215 26.885 275.785 ;
  END
 END i50
 PIN i51
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 267.045 26.885 267.615 ;
  END
 END i51
 PIN i52
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 240.635 26.885 241.205 ;
  END
 END i52
 PIN i53
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 285.095 26.885 285.665 ;
  END
 END i53
 PIN i54
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 281.105 27.645 281.675 ;
  END
 END i54
 PIN i55
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 276.925 26.885 277.495 ;
  END
 END i55
 PIN i56
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 297.445 27.645 298.015 ;
  END
 END i56
 PIN i57
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 293.265 26.885 293.835 ;
  END
 END i57
 PIN i58
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 217.835 26.885 218.405 ;
  END
 END i58
 PIN i59
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 213.845 27.645 214.415 ;
  END
 END i59
 PIN i60
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 209.665 26.885 210.235 ;
  END
 END i60
 PIN i61
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 205.675 27.645 206.245 ;
  END
 END i61
 PIN i62
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 226.005 26.885 226.575 ;
  END
 END i62
 PIN i63
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 109.155 26.885 109.725 ;
  END
 END i63
 PIN i64
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 113.145 27.645 113.715 ;
  END
 END i64
 PIN i65
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 117.325 26.885 117.895 ;
  END
 END i65
 PIN i66
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 121.315 27.645 121.885 ;
  END
 END i66
 PIN i67
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 100.985 26.885 101.555 ;
  END
 END i67
 PIN i68
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 41.895 26.885 42.465 ;
  END
 END i68
 PIN i69
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 45.885 27.645 46.455 ;
  END
 END i69
 PIN i70
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 50.065 26.885 50.635 ;
  END
 END i70
 PIN i71
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 33.725 26.885 34.295 ;
  END
 END i71
 PIN i72
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 54.055 27.645 54.625 ;
  END
 END i72
 PIN i73
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 289.275 27.645 289.845 ;
  END
 END i73
 PIN i74
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 222.015 27.645 222.585 ;
  END
 END i74
 PIN i75
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 104.975 27.645 105.545 ;
  END
 END i75
 PIN i76
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 37.715 27.645 38.285 ;
  END
 END i76
 PIN i77
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 18.335 175.845 18.905 176.415 ;
  END
 END i77
 PIN i78
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 18.335 162.545 18.905 163.115 ;
  END
 END i78
 PIN i79
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 331.835 27.645 332.405 ;
  END
 END i79
 PIN i80
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 323.665 27.645 324.235 ;
  END
 END i80
 PIN i81
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 231.895 27.645 232.465 ;
  END
 END i81
 PIN i82
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 223.725 27.645 224.295 ;
  END
 END i82
 PIN i83
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 215.555 27.645 216.125 ;
  END
 END i83
 PIN i84
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 207.385 27.645 207.955 ;
  END
 END i84
 PIN i85
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 199.215 27.645 199.785 ;
  END
 END i85
 PIN i86
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 191.045 27.645 191.615 ;
  END
 END i86
 PIN i87
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 182.875 27.645 183.445 ;
  END
 END i87
 PIN i88
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 144.115 27.645 144.685 ;
  END
 END i88
 PIN i89
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 135.945 27.645 136.515 ;
  END
 END i89
 PIN i90
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 127.775 27.645 128.345 ;
  END
 END i90
 PIN i91
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 315.495 27.645 316.065 ;
  END
 END i91
 PIN i92
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 119.605 27.645 120.175 ;
  END
 END i92
 PIN i93
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 111.435 27.645 112.005 ;
  END
 END i93
 PIN i94
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 103.265 27.645 103.835 ;
  END
 END i94
 PIN i95
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 95.095 27.645 95.665 ;
  END
 END i95
 PIN i96
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 86.925 27.645 87.495 ;
  END
 END i96
 PIN i97
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 60.515 27.645 61.085 ;
  END
 END i97
 PIN i98
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 52.345 27.645 52.915 ;
  END
 END i98
 PIN i99
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 44.175 27.645 44.745 ;
  END
 END i99
 PIN i100
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 36.005 27.645 36.575 ;
  END
 END i100
 PIN i101
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 27.835 27.645 28.405 ;
  END
 END i101
 PIN i102
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 307.325 27.645 307.895 ;
  END
 END i102
 PIN i103
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 19.665 27.645 20.235 ;
  END
 END i103
 PIN i104
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 11.495 27.645 12.065 ;
  END
 END i104
 PIN i105
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 3.325 27.645 3.895 ;
  END
 END i105
 PIN i106
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 299.155 27.645 299.725 ;
  END
 END i106
 PIN i107
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 290.985 27.645 291.555 ;
  END
 END i107
 PIN i108
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 282.815 27.645 283.385 ;
  END
 END i108
 PIN i109
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 274.645 27.645 275.215 ;
  END
 END i109
 PIN i110
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 266.475 27.645 267.045 ;
  END
 END i110
 PIN i111
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 240.065 27.645 240.635 ;
  END
 END i111
 PIN i112
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 168.245 3.705 168.815 ;
  END
 END i112
 PIN i113
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 167.865 4.465 168.435 ;
  END
 END i113
 PIN i114
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 331.265 28.405 331.835 ;
  END
 END i114
 PIN i115
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 323.095 28.405 323.665 ;
  END
 END i115
 PIN i116
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 231.325 28.405 231.895 ;
  END
 END i116
 PIN i117
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 223.155 28.405 223.725 ;
  END
 END i117
 PIN i118
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 214.985 28.405 215.555 ;
  END
 END i118
 PIN i119
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 206.815 28.405 207.385 ;
  END
 END i119
 PIN i120
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 198.645 28.405 199.215 ;
  END
 END i120
 PIN i121
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 190.475 28.405 191.045 ;
  END
 END i121
 PIN i122
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 182.305 28.405 182.875 ;
  END
 END i122
 PIN i123
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 144.685 28.405 145.255 ;
  END
 END i123
 PIN i124
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 136.515 28.405 137.085 ;
  END
 END i124
 PIN i125
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 128.345 28.405 128.915 ;
  END
 END i125
 PIN i126
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 314.925 28.405 315.495 ;
  END
 END i126
 PIN i127
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 120.175 28.405 120.745 ;
  END
 END i127
 PIN i128
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 112.005 28.405 112.575 ;
  END
 END i128
 PIN i129
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 103.835 28.405 104.405 ;
  END
 END i129
 PIN i130
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 95.665 28.405 96.235 ;
  END
 END i130
 PIN i131
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 87.495 28.405 88.065 ;
  END
 END i131
 PIN i132
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 61.085 28.405 61.655 ;
  END
 END i132
 PIN i133
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 52.915 28.405 53.485 ;
  END
 END i133
 PIN i134
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 44.745 28.405 45.315 ;
  END
 END i134
 PIN i135
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 36.575 28.405 37.145 ;
  END
 END i135
 PIN i136
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 28.405 28.405 28.975 ;
  END
 END i136
 PIN i137
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 306.755 28.405 307.325 ;
  END
 END i137
 PIN i138
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 20.235 28.405 20.805 ;
  END
 END i138
 PIN i139
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 12.065 28.405 12.635 ;
  END
 END i139
 PIN i140
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 3.895 28.405 4.465 ;
  END
 END i140
 PIN i141
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 298.585 28.405 299.155 ;
  END
 END i141
 PIN i142
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 290.415 28.405 290.985 ;
  END
 END i142
 PIN i143
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 282.245 28.405 282.815 ;
  END
 END i143
 PIN i144
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 274.075 28.405 274.645 ;
  END
 END i144
 PIN i145
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 265.905 28.405 266.475 ;
  END
 END i145
 PIN i146
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 239.495 28.405 240.065 ;
  END
 END i146
 PIN i147
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 4.275 175.845 4.845 176.415 ;
  END
 END i147
 PIN i148
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 5.415 175.845 5.985 176.415 ;
  END
 END i148
 PIN i149
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 7.315 175.845 7.885 176.415 ;
  END
 END i149
 PIN i150
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 8.835 175.845 9.405 176.415 ;
  END
 END i150
 PIN i151
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 175.845 10.925 176.415 ;
  END
 END i151
 PIN i152
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 11.875 175.845 12.445 176.415 ;
  END
 END i152
 PIN i153
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 4.275 162.545 4.845 163.115 ;
  END
 END i153
 PIN i154
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 5.415 162.545 5.985 163.115 ;
  END
 END i154
 PIN i155
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 7.315 162.545 7.885 163.115 ;
  END
 END i155
 PIN i156
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 8.835 162.545 9.405 163.115 ;
  END
 END i156
 PIN i157
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 162.545 10.925 163.115 ;
  END
 END i157
 PIN i158
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 11.875 162.545 12.445 163.115 ;
  END
 END i158
 OBS
  LAYER metal1 ;
   RECT 23.18 0.0 508.44 1.71 ;
   RECT 23.18 1.71 508.44 3.42 ;
   RECT 23.18 3.42 508.44 5.13 ;
   RECT 23.18 5.13 508.44 6.84 ;
   RECT 23.18 6.84 508.44 8.55 ;
   RECT 23.18 8.55 508.44 10.26 ;
   RECT 23.18 10.26 508.44 11.97 ;
   RECT 23.18 11.97 508.44 13.68 ;
   RECT 23.18 13.68 508.44 15.39 ;
   RECT 23.18 15.39 508.44 17.1 ;
   RECT 23.18 17.1 508.44 18.81 ;
   RECT 23.18 18.81 508.44 20.52 ;
   RECT 23.18 20.52 508.44 22.23 ;
   RECT 23.18 22.23 508.44 23.94 ;
   RECT 23.18 23.94 508.44 25.65 ;
   RECT 23.18 25.65 508.44 27.36 ;
   RECT 23.18 27.36 508.44 29.07 ;
   RECT 23.18 29.07 508.44 30.78 ;
   RECT 23.18 30.78 508.44 32.49 ;
   RECT 23.18 32.49 508.44 34.2 ;
   RECT 23.18 34.2 508.44 35.91 ;
   RECT 23.18 35.91 508.44 37.62 ;
   RECT 23.18 37.62 508.44 39.33 ;
   RECT 23.18 39.33 508.44 41.04 ;
   RECT 23.18 41.04 508.44 42.75 ;
   RECT 23.18 42.75 508.44 44.46 ;
   RECT 23.18 44.46 508.44 46.17 ;
   RECT 23.18 46.17 508.44 47.88 ;
   RECT 23.18 47.88 508.44 49.59 ;
   RECT 23.18 49.59 508.44 51.3 ;
   RECT 23.18 51.3 508.44 53.01 ;
   RECT 23.18 53.01 508.44 54.72 ;
   RECT 23.18 54.72 508.44 56.43 ;
   RECT 23.18 56.43 508.44 58.14 ;
   RECT 23.18 58.14 508.44 59.85 ;
   RECT 23.18 59.85 508.44 61.56 ;
   RECT 23.18 61.56 508.44 63.27 ;
   RECT 23.18 63.27 508.44 64.98 ;
   RECT 23.18 64.98 508.44 66.69 ;
   RECT 23.18 66.69 508.44 68.4 ;
   RECT 23.18 68.4 508.44 70.11 ;
   RECT 23.18 70.11 508.44 71.82 ;
   RECT 23.18 71.82 508.44 73.53 ;
   RECT 23.18 73.53 508.44 75.24 ;
   RECT 23.18 75.24 508.44 76.95 ;
   RECT 23.18 76.95 508.44 78.66 ;
   RECT 23.18 78.66 508.44 80.37 ;
   RECT 23.18 80.37 508.44 82.08 ;
   RECT 23.18 82.08 508.44 83.79 ;
   RECT 23.18 83.79 508.44 85.5 ;
   RECT 23.18 85.5 508.44 87.21 ;
   RECT 23.18 87.21 508.44 88.92 ;
   RECT 23.18 88.92 508.44 90.63 ;
   RECT 23.18 90.63 508.44 92.34 ;
   RECT 23.18 92.34 508.44 94.05 ;
   RECT 23.18 94.05 508.44 95.76 ;
   RECT 23.18 95.76 508.44 97.47 ;
   RECT 23.18 97.47 508.44 99.18 ;
   RECT 23.18 99.18 508.44 100.89 ;
   RECT 23.18 100.89 508.44 102.6 ;
   RECT 23.18 102.6 508.44 104.31 ;
   RECT 23.18 104.31 508.44 106.02 ;
   RECT 23.18 106.02 508.44 107.73 ;
   RECT 23.18 107.73 508.44 109.44 ;
   RECT 23.18 109.44 508.44 111.15 ;
   RECT 23.18 111.15 508.44 112.86 ;
   RECT 23.18 112.86 508.44 114.57 ;
   RECT 23.18 114.57 508.44 116.28 ;
   RECT 23.18 116.28 508.44 117.99 ;
   RECT 23.18 117.99 508.44 119.7 ;
   RECT 23.18 119.7 508.44 121.41 ;
   RECT 23.18 121.41 508.44 123.12 ;
   RECT 23.18 123.12 508.44 124.83 ;
   RECT 23.18 124.83 508.44 126.54 ;
   RECT 23.18 126.54 508.44 128.25 ;
   RECT 23.18 128.25 508.44 129.96 ;
   RECT 23.18 129.96 508.44 131.67 ;
   RECT 23.18 131.67 508.44 133.38 ;
   RECT 23.18 133.38 508.44 135.09 ;
   RECT 23.18 135.09 508.44 136.8 ;
   RECT 23.18 136.8 508.44 138.51 ;
   RECT 23.18 138.51 508.44 140.22 ;
   RECT 23.18 140.22 508.44 141.93 ;
   RECT 23.18 141.93 508.44 143.64 ;
   RECT 23.18 143.64 508.44 145.35 ;
   RECT 23.18 145.35 508.44 147.06 ;
   RECT 23.18 147.06 508.44 148.77 ;
   RECT 23.18 148.77 508.44 150.48 ;
   RECT 0.0 150.48 508.44 152.19 ;
   RECT 0.0 152.19 508.44 153.9 ;
   RECT 0.0 153.9 508.44 155.61 ;
   RECT 0.0 155.61 508.44 157.32 ;
   RECT 0.0 157.32 508.44 159.03 ;
   RECT 0.0 159.03 508.44 160.74 ;
   RECT 0.0 160.74 508.44 162.45 ;
   RECT 0.0 162.45 508.44 164.16 ;
   RECT 0.0 164.16 508.44 165.87 ;
   RECT 0.0 165.87 508.44 167.58 ;
   RECT 0.0 167.58 508.44 169.29 ;
   RECT 0.0 169.29 508.44 171.0 ;
   RECT 0.0 171.0 508.44 172.71 ;
   RECT 0.0 172.71 508.44 174.42 ;
   RECT 0.0 174.42 508.44 176.13 ;
   RECT 0.0 176.13 508.44 177.84 ;
   RECT 0.0 177.84 508.44 179.55 ;
   RECT 23.18 179.55 508.44 181.26 ;
   RECT 23.18 181.26 508.44 182.97 ;
   RECT 23.18 182.97 508.44 184.68 ;
   RECT 23.18 184.68 508.44 186.39 ;
   RECT 23.18 186.39 508.44 188.1 ;
   RECT 23.18 188.1 508.44 189.81 ;
   RECT 23.18 189.81 508.44 191.52 ;
   RECT 23.18 191.52 508.44 193.23 ;
   RECT 23.18 193.23 508.44 194.94 ;
   RECT 23.18 194.94 508.44 196.65 ;
   RECT 23.18 196.65 508.44 198.36 ;
   RECT 23.18 198.36 508.44 200.07 ;
   RECT 23.18 200.07 508.44 201.78 ;
   RECT 23.18 201.78 508.44 203.49 ;
   RECT 23.18 203.49 508.44 205.2 ;
   RECT 23.18 205.2 508.44 206.91 ;
   RECT 23.18 206.91 508.44 208.62 ;
   RECT 23.18 208.62 508.44 210.33 ;
   RECT 23.18 210.33 508.44 212.04 ;
   RECT 23.18 212.04 508.44 213.75 ;
   RECT 23.18 213.75 508.44 215.46 ;
   RECT 23.18 215.46 508.44 217.17 ;
   RECT 23.18 217.17 508.44 218.88 ;
   RECT 23.18 218.88 508.44 220.59 ;
   RECT 23.18 220.59 508.44 222.3 ;
   RECT 23.18 222.3 508.44 224.01 ;
   RECT 23.18 224.01 508.44 225.72 ;
   RECT 23.18 225.72 508.44 227.43 ;
   RECT 23.18 227.43 508.44 229.14 ;
   RECT 23.18 229.14 508.44 230.85 ;
   RECT 23.18 230.85 508.44 232.56 ;
   RECT 23.18 232.56 508.44 234.27 ;
   RECT 23.18 234.27 508.44 235.98 ;
   RECT 23.18 235.98 508.44 237.69 ;
   RECT 23.18 237.69 508.44 239.4 ;
   RECT 23.18 239.4 508.44 241.11 ;
   RECT 23.18 241.11 508.44 242.82 ;
   RECT 23.18 242.82 508.44 244.53 ;
   RECT 23.18 244.53 508.44 246.24 ;
   RECT 23.18 246.24 508.44 247.95 ;
   RECT 23.18 247.95 508.44 249.66 ;
   RECT 23.18 249.66 508.44 251.37 ;
   RECT 23.18 251.37 508.44 253.08 ;
   RECT 23.18 253.08 508.44 254.79 ;
   RECT 23.18 254.79 508.44 256.5 ;
   RECT 23.18 256.5 508.44 258.21 ;
   RECT 23.18 258.21 508.44 259.92 ;
   RECT 23.18 259.92 508.44 261.63 ;
   RECT 23.18 261.63 508.44 263.34 ;
   RECT 23.18 263.34 508.44 265.05 ;
   RECT 23.18 265.05 508.44 266.76 ;
   RECT 23.18 266.76 508.44 268.47 ;
   RECT 23.18 268.47 508.44 270.18 ;
   RECT 23.18 270.18 508.44 271.89 ;
   RECT 23.18 271.89 508.44 273.6 ;
   RECT 23.18 273.6 508.44 275.31 ;
   RECT 23.18 275.31 508.44 277.02 ;
   RECT 23.18 277.02 508.44 278.73 ;
   RECT 23.18 278.73 508.44 280.44 ;
   RECT 23.18 280.44 508.44 282.15 ;
   RECT 23.18 282.15 508.44 283.86 ;
   RECT 23.18 283.86 508.44 285.57 ;
   RECT 23.18 285.57 508.44 287.28 ;
   RECT 23.18 287.28 508.44 288.99 ;
   RECT 23.18 288.99 508.44 290.7 ;
   RECT 23.18 290.7 508.44 292.41 ;
   RECT 23.18 292.41 508.44 294.12 ;
   RECT 23.18 294.12 508.44 295.83 ;
   RECT 23.18 295.83 508.44 297.54 ;
   RECT 23.18 297.54 508.44 299.25 ;
   RECT 23.18 299.25 508.44 300.96 ;
   RECT 23.18 300.96 508.44 302.67 ;
   RECT 23.18 302.67 508.44 304.38 ;
   RECT 23.18 304.38 508.44 306.09 ;
   RECT 23.18 306.09 508.44 307.8 ;
   RECT 23.18 307.8 508.44 309.51 ;
   RECT 23.18 309.51 508.44 311.22 ;
   RECT 23.18 311.22 508.44 312.93 ;
   RECT 23.18 312.93 508.44 314.64 ;
   RECT 23.18 314.64 508.44 316.35 ;
   RECT 23.18 316.35 508.44 318.06 ;
   RECT 23.18 318.06 508.44 319.77 ;
   RECT 23.18 319.77 508.44 321.48 ;
   RECT 23.18 321.48 508.44 323.19 ;
   RECT 23.18 323.19 508.44 324.9 ;
   RECT 23.18 324.9 508.44 326.61 ;
   RECT 23.18 326.61 508.44 328.32 ;
   RECT 23.18 328.32 508.44 330.03 ;
   RECT 23.18 330.03 508.44 331.74 ;
   RECT 23.18 331.74 508.44 333.45 ;
   RECT 23.18 333.45 508.44 335.16 ;
   RECT 23.18 335.16 508.44 336.87 ;
  LAYER via1 ;
   RECT 23.18 0.0 508.44 1.71 ;
   RECT 23.18 1.71 508.44 3.42 ;
   RECT 23.18 3.42 508.44 5.13 ;
   RECT 23.18 5.13 508.44 6.84 ;
   RECT 23.18 6.84 508.44 8.55 ;
   RECT 23.18 8.55 508.44 10.26 ;
   RECT 23.18 10.26 508.44 11.97 ;
   RECT 23.18 11.97 508.44 13.68 ;
   RECT 23.18 13.68 508.44 15.39 ;
   RECT 23.18 15.39 508.44 17.1 ;
   RECT 23.18 17.1 508.44 18.81 ;
   RECT 23.18 18.81 508.44 20.52 ;
   RECT 23.18 20.52 508.44 22.23 ;
   RECT 23.18 22.23 508.44 23.94 ;
   RECT 23.18 23.94 508.44 25.65 ;
   RECT 23.18 25.65 508.44 27.36 ;
   RECT 23.18 27.36 508.44 29.07 ;
   RECT 23.18 29.07 508.44 30.78 ;
   RECT 23.18 30.78 508.44 32.49 ;
   RECT 23.18 32.49 508.44 34.2 ;
   RECT 23.18 34.2 508.44 35.91 ;
   RECT 23.18 35.91 508.44 37.62 ;
   RECT 23.18 37.62 508.44 39.33 ;
   RECT 23.18 39.33 508.44 41.04 ;
   RECT 23.18 41.04 508.44 42.75 ;
   RECT 23.18 42.75 508.44 44.46 ;
   RECT 23.18 44.46 508.44 46.17 ;
   RECT 23.18 46.17 508.44 47.88 ;
   RECT 23.18 47.88 508.44 49.59 ;
   RECT 23.18 49.59 508.44 51.3 ;
   RECT 23.18 51.3 508.44 53.01 ;
   RECT 23.18 53.01 508.44 54.72 ;
   RECT 23.18 54.72 508.44 56.43 ;
   RECT 23.18 56.43 508.44 58.14 ;
   RECT 23.18 58.14 508.44 59.85 ;
   RECT 23.18 59.85 508.44 61.56 ;
   RECT 23.18 61.56 508.44 63.27 ;
   RECT 23.18 63.27 508.44 64.98 ;
   RECT 23.18 64.98 508.44 66.69 ;
   RECT 23.18 66.69 508.44 68.4 ;
   RECT 23.18 68.4 508.44 70.11 ;
   RECT 23.18 70.11 508.44 71.82 ;
   RECT 23.18 71.82 508.44 73.53 ;
   RECT 23.18 73.53 508.44 75.24 ;
   RECT 23.18 75.24 508.44 76.95 ;
   RECT 23.18 76.95 508.44 78.66 ;
   RECT 23.18 78.66 508.44 80.37 ;
   RECT 23.18 80.37 508.44 82.08 ;
   RECT 23.18 82.08 508.44 83.79 ;
   RECT 23.18 83.79 508.44 85.5 ;
   RECT 23.18 85.5 508.44 87.21 ;
   RECT 23.18 87.21 508.44 88.92 ;
   RECT 23.18 88.92 508.44 90.63 ;
   RECT 23.18 90.63 508.44 92.34 ;
   RECT 23.18 92.34 508.44 94.05 ;
   RECT 23.18 94.05 508.44 95.76 ;
   RECT 23.18 95.76 508.44 97.47 ;
   RECT 23.18 97.47 508.44 99.18 ;
   RECT 23.18 99.18 508.44 100.89 ;
   RECT 23.18 100.89 508.44 102.6 ;
   RECT 23.18 102.6 508.44 104.31 ;
   RECT 23.18 104.31 508.44 106.02 ;
   RECT 23.18 106.02 508.44 107.73 ;
   RECT 23.18 107.73 508.44 109.44 ;
   RECT 23.18 109.44 508.44 111.15 ;
   RECT 23.18 111.15 508.44 112.86 ;
   RECT 23.18 112.86 508.44 114.57 ;
   RECT 23.18 114.57 508.44 116.28 ;
   RECT 23.18 116.28 508.44 117.99 ;
   RECT 23.18 117.99 508.44 119.7 ;
   RECT 23.18 119.7 508.44 121.41 ;
   RECT 23.18 121.41 508.44 123.12 ;
   RECT 23.18 123.12 508.44 124.83 ;
   RECT 23.18 124.83 508.44 126.54 ;
   RECT 23.18 126.54 508.44 128.25 ;
   RECT 23.18 128.25 508.44 129.96 ;
   RECT 23.18 129.96 508.44 131.67 ;
   RECT 23.18 131.67 508.44 133.38 ;
   RECT 23.18 133.38 508.44 135.09 ;
   RECT 23.18 135.09 508.44 136.8 ;
   RECT 23.18 136.8 508.44 138.51 ;
   RECT 23.18 138.51 508.44 140.22 ;
   RECT 23.18 140.22 508.44 141.93 ;
   RECT 23.18 141.93 508.44 143.64 ;
   RECT 23.18 143.64 508.44 145.35 ;
   RECT 23.18 145.35 508.44 147.06 ;
   RECT 23.18 147.06 508.44 148.77 ;
   RECT 23.18 148.77 508.44 150.48 ;
   RECT 0.0 150.48 508.44 152.19 ;
   RECT 0.0 152.19 508.44 153.9 ;
   RECT 0.0 153.9 508.44 155.61 ;
   RECT 0.0 155.61 508.44 157.32 ;
   RECT 0.0 157.32 508.44 159.03 ;
   RECT 0.0 159.03 508.44 160.74 ;
   RECT 0.0 160.74 508.44 162.45 ;
   RECT 0.0 162.45 508.44 164.16 ;
   RECT 0.0 164.16 508.44 165.87 ;
   RECT 0.0 165.87 508.44 167.58 ;
   RECT 0.0 167.58 508.44 169.29 ;
   RECT 0.0 169.29 508.44 171.0 ;
   RECT 0.0 171.0 508.44 172.71 ;
   RECT 0.0 172.71 508.44 174.42 ;
   RECT 0.0 174.42 508.44 176.13 ;
   RECT 0.0 176.13 508.44 177.84 ;
   RECT 0.0 177.84 508.44 179.55 ;
   RECT 23.18 179.55 508.44 181.26 ;
   RECT 23.18 181.26 508.44 182.97 ;
   RECT 23.18 182.97 508.44 184.68 ;
   RECT 23.18 184.68 508.44 186.39 ;
   RECT 23.18 186.39 508.44 188.1 ;
   RECT 23.18 188.1 508.44 189.81 ;
   RECT 23.18 189.81 508.44 191.52 ;
   RECT 23.18 191.52 508.44 193.23 ;
   RECT 23.18 193.23 508.44 194.94 ;
   RECT 23.18 194.94 508.44 196.65 ;
   RECT 23.18 196.65 508.44 198.36 ;
   RECT 23.18 198.36 508.44 200.07 ;
   RECT 23.18 200.07 508.44 201.78 ;
   RECT 23.18 201.78 508.44 203.49 ;
   RECT 23.18 203.49 508.44 205.2 ;
   RECT 23.18 205.2 508.44 206.91 ;
   RECT 23.18 206.91 508.44 208.62 ;
   RECT 23.18 208.62 508.44 210.33 ;
   RECT 23.18 210.33 508.44 212.04 ;
   RECT 23.18 212.04 508.44 213.75 ;
   RECT 23.18 213.75 508.44 215.46 ;
   RECT 23.18 215.46 508.44 217.17 ;
   RECT 23.18 217.17 508.44 218.88 ;
   RECT 23.18 218.88 508.44 220.59 ;
   RECT 23.18 220.59 508.44 222.3 ;
   RECT 23.18 222.3 508.44 224.01 ;
   RECT 23.18 224.01 508.44 225.72 ;
   RECT 23.18 225.72 508.44 227.43 ;
   RECT 23.18 227.43 508.44 229.14 ;
   RECT 23.18 229.14 508.44 230.85 ;
   RECT 23.18 230.85 508.44 232.56 ;
   RECT 23.18 232.56 508.44 234.27 ;
   RECT 23.18 234.27 508.44 235.98 ;
   RECT 23.18 235.98 508.44 237.69 ;
   RECT 23.18 237.69 508.44 239.4 ;
   RECT 23.18 239.4 508.44 241.11 ;
   RECT 23.18 241.11 508.44 242.82 ;
   RECT 23.18 242.82 508.44 244.53 ;
   RECT 23.18 244.53 508.44 246.24 ;
   RECT 23.18 246.24 508.44 247.95 ;
   RECT 23.18 247.95 508.44 249.66 ;
   RECT 23.18 249.66 508.44 251.37 ;
   RECT 23.18 251.37 508.44 253.08 ;
   RECT 23.18 253.08 508.44 254.79 ;
   RECT 23.18 254.79 508.44 256.5 ;
   RECT 23.18 256.5 508.44 258.21 ;
   RECT 23.18 258.21 508.44 259.92 ;
   RECT 23.18 259.92 508.44 261.63 ;
   RECT 23.18 261.63 508.44 263.34 ;
   RECT 23.18 263.34 508.44 265.05 ;
   RECT 23.18 265.05 508.44 266.76 ;
   RECT 23.18 266.76 508.44 268.47 ;
   RECT 23.18 268.47 508.44 270.18 ;
   RECT 23.18 270.18 508.44 271.89 ;
   RECT 23.18 271.89 508.44 273.6 ;
   RECT 23.18 273.6 508.44 275.31 ;
   RECT 23.18 275.31 508.44 277.02 ;
   RECT 23.18 277.02 508.44 278.73 ;
   RECT 23.18 278.73 508.44 280.44 ;
   RECT 23.18 280.44 508.44 282.15 ;
   RECT 23.18 282.15 508.44 283.86 ;
   RECT 23.18 283.86 508.44 285.57 ;
   RECT 23.18 285.57 508.44 287.28 ;
   RECT 23.18 287.28 508.44 288.99 ;
   RECT 23.18 288.99 508.44 290.7 ;
   RECT 23.18 290.7 508.44 292.41 ;
   RECT 23.18 292.41 508.44 294.12 ;
   RECT 23.18 294.12 508.44 295.83 ;
   RECT 23.18 295.83 508.44 297.54 ;
   RECT 23.18 297.54 508.44 299.25 ;
   RECT 23.18 299.25 508.44 300.96 ;
   RECT 23.18 300.96 508.44 302.67 ;
   RECT 23.18 302.67 508.44 304.38 ;
   RECT 23.18 304.38 508.44 306.09 ;
   RECT 23.18 306.09 508.44 307.8 ;
   RECT 23.18 307.8 508.44 309.51 ;
   RECT 23.18 309.51 508.44 311.22 ;
   RECT 23.18 311.22 508.44 312.93 ;
   RECT 23.18 312.93 508.44 314.64 ;
   RECT 23.18 314.64 508.44 316.35 ;
   RECT 23.18 316.35 508.44 318.06 ;
   RECT 23.18 318.06 508.44 319.77 ;
   RECT 23.18 319.77 508.44 321.48 ;
   RECT 23.18 321.48 508.44 323.19 ;
   RECT 23.18 323.19 508.44 324.9 ;
   RECT 23.18 324.9 508.44 326.61 ;
   RECT 23.18 326.61 508.44 328.32 ;
   RECT 23.18 328.32 508.44 330.03 ;
   RECT 23.18 330.03 508.44 331.74 ;
   RECT 23.18 331.74 508.44 333.45 ;
   RECT 23.18 333.45 508.44 335.16 ;
   RECT 23.18 335.16 508.44 336.87 ;
  LAYER metal2 ;
   RECT 23.18 0.0 508.44 1.71 ;
   RECT 23.18 1.71 508.44 3.42 ;
   RECT 23.18 3.42 508.44 5.13 ;
   RECT 23.18 5.13 508.44 6.84 ;
   RECT 23.18 6.84 508.44 8.55 ;
   RECT 23.18 8.55 508.44 10.26 ;
   RECT 23.18 10.26 508.44 11.97 ;
   RECT 23.18 11.97 508.44 13.68 ;
   RECT 23.18 13.68 508.44 15.39 ;
   RECT 23.18 15.39 508.44 17.1 ;
   RECT 23.18 17.1 508.44 18.81 ;
   RECT 23.18 18.81 508.44 20.52 ;
   RECT 23.18 20.52 508.44 22.23 ;
   RECT 23.18 22.23 508.44 23.94 ;
   RECT 23.18 23.94 508.44 25.65 ;
   RECT 23.18 25.65 508.44 27.36 ;
   RECT 23.18 27.36 508.44 29.07 ;
   RECT 23.18 29.07 508.44 30.78 ;
   RECT 23.18 30.78 508.44 32.49 ;
   RECT 23.18 32.49 508.44 34.2 ;
   RECT 23.18 34.2 508.44 35.91 ;
   RECT 23.18 35.91 508.44 37.62 ;
   RECT 23.18 37.62 508.44 39.33 ;
   RECT 23.18 39.33 508.44 41.04 ;
   RECT 23.18 41.04 508.44 42.75 ;
   RECT 23.18 42.75 508.44 44.46 ;
   RECT 23.18 44.46 508.44 46.17 ;
   RECT 23.18 46.17 508.44 47.88 ;
   RECT 23.18 47.88 508.44 49.59 ;
   RECT 23.18 49.59 508.44 51.3 ;
   RECT 23.18 51.3 508.44 53.01 ;
   RECT 23.18 53.01 508.44 54.72 ;
   RECT 23.18 54.72 508.44 56.43 ;
   RECT 23.18 56.43 508.44 58.14 ;
   RECT 23.18 58.14 508.44 59.85 ;
   RECT 23.18 59.85 508.44 61.56 ;
   RECT 23.18 61.56 508.44 63.27 ;
   RECT 23.18 63.27 508.44 64.98 ;
   RECT 23.18 64.98 508.44 66.69 ;
   RECT 23.18 66.69 508.44 68.4 ;
   RECT 23.18 68.4 508.44 70.11 ;
   RECT 23.18 70.11 508.44 71.82 ;
   RECT 23.18 71.82 508.44 73.53 ;
   RECT 23.18 73.53 508.44 75.24 ;
   RECT 23.18 75.24 508.44 76.95 ;
   RECT 23.18 76.95 508.44 78.66 ;
   RECT 23.18 78.66 508.44 80.37 ;
   RECT 23.18 80.37 508.44 82.08 ;
   RECT 23.18 82.08 508.44 83.79 ;
   RECT 23.18 83.79 508.44 85.5 ;
   RECT 23.18 85.5 508.44 87.21 ;
   RECT 23.18 87.21 508.44 88.92 ;
   RECT 23.18 88.92 508.44 90.63 ;
   RECT 23.18 90.63 508.44 92.34 ;
   RECT 23.18 92.34 508.44 94.05 ;
   RECT 23.18 94.05 508.44 95.76 ;
   RECT 23.18 95.76 508.44 97.47 ;
   RECT 23.18 97.47 508.44 99.18 ;
   RECT 23.18 99.18 508.44 100.89 ;
   RECT 23.18 100.89 508.44 102.6 ;
   RECT 23.18 102.6 508.44 104.31 ;
   RECT 23.18 104.31 508.44 106.02 ;
   RECT 23.18 106.02 508.44 107.73 ;
   RECT 23.18 107.73 508.44 109.44 ;
   RECT 23.18 109.44 508.44 111.15 ;
   RECT 23.18 111.15 508.44 112.86 ;
   RECT 23.18 112.86 508.44 114.57 ;
   RECT 23.18 114.57 508.44 116.28 ;
   RECT 23.18 116.28 508.44 117.99 ;
   RECT 23.18 117.99 508.44 119.7 ;
   RECT 23.18 119.7 508.44 121.41 ;
   RECT 23.18 121.41 508.44 123.12 ;
   RECT 23.18 123.12 508.44 124.83 ;
   RECT 23.18 124.83 508.44 126.54 ;
   RECT 23.18 126.54 508.44 128.25 ;
   RECT 23.18 128.25 508.44 129.96 ;
   RECT 23.18 129.96 508.44 131.67 ;
   RECT 23.18 131.67 508.44 133.38 ;
   RECT 23.18 133.38 508.44 135.09 ;
   RECT 23.18 135.09 508.44 136.8 ;
   RECT 23.18 136.8 508.44 138.51 ;
   RECT 23.18 138.51 508.44 140.22 ;
   RECT 23.18 140.22 508.44 141.93 ;
   RECT 23.18 141.93 508.44 143.64 ;
   RECT 23.18 143.64 508.44 145.35 ;
   RECT 23.18 145.35 508.44 147.06 ;
   RECT 23.18 147.06 508.44 148.77 ;
   RECT 23.18 148.77 508.44 150.48 ;
   RECT 0.0 150.48 508.44 152.19 ;
   RECT 0.0 152.19 508.44 153.9 ;
   RECT 0.0 153.9 508.44 155.61 ;
   RECT 0.0 155.61 508.44 157.32 ;
   RECT 0.0 157.32 508.44 159.03 ;
   RECT 0.0 159.03 508.44 160.74 ;
   RECT 0.0 160.74 508.44 162.45 ;
   RECT 0.0 162.45 508.44 164.16 ;
   RECT 0.0 164.16 508.44 165.87 ;
   RECT 0.0 165.87 508.44 167.58 ;
   RECT 0.0 167.58 508.44 169.29 ;
   RECT 0.0 169.29 508.44 171.0 ;
   RECT 0.0 171.0 508.44 172.71 ;
   RECT 0.0 172.71 508.44 174.42 ;
   RECT 0.0 174.42 508.44 176.13 ;
   RECT 0.0 176.13 508.44 177.84 ;
   RECT 0.0 177.84 508.44 179.55 ;
   RECT 23.18 179.55 508.44 181.26 ;
   RECT 23.18 181.26 508.44 182.97 ;
   RECT 23.18 182.97 508.44 184.68 ;
   RECT 23.18 184.68 508.44 186.39 ;
   RECT 23.18 186.39 508.44 188.1 ;
   RECT 23.18 188.1 508.44 189.81 ;
   RECT 23.18 189.81 508.44 191.52 ;
   RECT 23.18 191.52 508.44 193.23 ;
   RECT 23.18 193.23 508.44 194.94 ;
   RECT 23.18 194.94 508.44 196.65 ;
   RECT 23.18 196.65 508.44 198.36 ;
   RECT 23.18 198.36 508.44 200.07 ;
   RECT 23.18 200.07 508.44 201.78 ;
   RECT 23.18 201.78 508.44 203.49 ;
   RECT 23.18 203.49 508.44 205.2 ;
   RECT 23.18 205.2 508.44 206.91 ;
   RECT 23.18 206.91 508.44 208.62 ;
   RECT 23.18 208.62 508.44 210.33 ;
   RECT 23.18 210.33 508.44 212.04 ;
   RECT 23.18 212.04 508.44 213.75 ;
   RECT 23.18 213.75 508.44 215.46 ;
   RECT 23.18 215.46 508.44 217.17 ;
   RECT 23.18 217.17 508.44 218.88 ;
   RECT 23.18 218.88 508.44 220.59 ;
   RECT 23.18 220.59 508.44 222.3 ;
   RECT 23.18 222.3 508.44 224.01 ;
   RECT 23.18 224.01 508.44 225.72 ;
   RECT 23.18 225.72 508.44 227.43 ;
   RECT 23.18 227.43 508.44 229.14 ;
   RECT 23.18 229.14 508.44 230.85 ;
   RECT 23.18 230.85 508.44 232.56 ;
   RECT 23.18 232.56 508.44 234.27 ;
   RECT 23.18 234.27 508.44 235.98 ;
   RECT 23.18 235.98 508.44 237.69 ;
   RECT 23.18 237.69 508.44 239.4 ;
   RECT 23.18 239.4 508.44 241.11 ;
   RECT 23.18 241.11 508.44 242.82 ;
   RECT 23.18 242.82 508.44 244.53 ;
   RECT 23.18 244.53 508.44 246.24 ;
   RECT 23.18 246.24 508.44 247.95 ;
   RECT 23.18 247.95 508.44 249.66 ;
   RECT 23.18 249.66 508.44 251.37 ;
   RECT 23.18 251.37 508.44 253.08 ;
   RECT 23.18 253.08 508.44 254.79 ;
   RECT 23.18 254.79 508.44 256.5 ;
   RECT 23.18 256.5 508.44 258.21 ;
   RECT 23.18 258.21 508.44 259.92 ;
   RECT 23.18 259.92 508.44 261.63 ;
   RECT 23.18 261.63 508.44 263.34 ;
   RECT 23.18 263.34 508.44 265.05 ;
   RECT 23.18 265.05 508.44 266.76 ;
   RECT 23.18 266.76 508.44 268.47 ;
   RECT 23.18 268.47 508.44 270.18 ;
   RECT 23.18 270.18 508.44 271.89 ;
   RECT 23.18 271.89 508.44 273.6 ;
   RECT 23.18 273.6 508.44 275.31 ;
   RECT 23.18 275.31 508.44 277.02 ;
   RECT 23.18 277.02 508.44 278.73 ;
   RECT 23.18 278.73 508.44 280.44 ;
   RECT 23.18 280.44 508.44 282.15 ;
   RECT 23.18 282.15 508.44 283.86 ;
   RECT 23.18 283.86 508.44 285.57 ;
   RECT 23.18 285.57 508.44 287.28 ;
   RECT 23.18 287.28 508.44 288.99 ;
   RECT 23.18 288.99 508.44 290.7 ;
   RECT 23.18 290.7 508.44 292.41 ;
   RECT 23.18 292.41 508.44 294.12 ;
   RECT 23.18 294.12 508.44 295.83 ;
   RECT 23.18 295.83 508.44 297.54 ;
   RECT 23.18 297.54 508.44 299.25 ;
   RECT 23.18 299.25 508.44 300.96 ;
   RECT 23.18 300.96 508.44 302.67 ;
   RECT 23.18 302.67 508.44 304.38 ;
   RECT 23.18 304.38 508.44 306.09 ;
   RECT 23.18 306.09 508.44 307.8 ;
   RECT 23.18 307.8 508.44 309.51 ;
   RECT 23.18 309.51 508.44 311.22 ;
   RECT 23.18 311.22 508.44 312.93 ;
   RECT 23.18 312.93 508.44 314.64 ;
   RECT 23.18 314.64 508.44 316.35 ;
   RECT 23.18 316.35 508.44 318.06 ;
   RECT 23.18 318.06 508.44 319.77 ;
   RECT 23.18 319.77 508.44 321.48 ;
   RECT 23.18 321.48 508.44 323.19 ;
   RECT 23.18 323.19 508.44 324.9 ;
   RECT 23.18 324.9 508.44 326.61 ;
   RECT 23.18 326.61 508.44 328.32 ;
   RECT 23.18 328.32 508.44 330.03 ;
   RECT 23.18 330.03 508.44 331.74 ;
   RECT 23.18 331.74 508.44 333.45 ;
   RECT 23.18 333.45 508.44 335.16 ;
   RECT 23.18 335.16 508.44 336.87 ;
  LAYER via2 ;
   RECT 23.18 0.0 508.44 1.71 ;
   RECT 23.18 1.71 508.44 3.42 ;
   RECT 23.18 3.42 508.44 5.13 ;
   RECT 23.18 5.13 508.44 6.84 ;
   RECT 23.18 6.84 508.44 8.55 ;
   RECT 23.18 8.55 508.44 10.26 ;
   RECT 23.18 10.26 508.44 11.97 ;
   RECT 23.18 11.97 508.44 13.68 ;
   RECT 23.18 13.68 508.44 15.39 ;
   RECT 23.18 15.39 508.44 17.1 ;
   RECT 23.18 17.1 508.44 18.81 ;
   RECT 23.18 18.81 508.44 20.52 ;
   RECT 23.18 20.52 508.44 22.23 ;
   RECT 23.18 22.23 508.44 23.94 ;
   RECT 23.18 23.94 508.44 25.65 ;
   RECT 23.18 25.65 508.44 27.36 ;
   RECT 23.18 27.36 508.44 29.07 ;
   RECT 23.18 29.07 508.44 30.78 ;
   RECT 23.18 30.78 508.44 32.49 ;
   RECT 23.18 32.49 508.44 34.2 ;
   RECT 23.18 34.2 508.44 35.91 ;
   RECT 23.18 35.91 508.44 37.62 ;
   RECT 23.18 37.62 508.44 39.33 ;
   RECT 23.18 39.33 508.44 41.04 ;
   RECT 23.18 41.04 508.44 42.75 ;
   RECT 23.18 42.75 508.44 44.46 ;
   RECT 23.18 44.46 508.44 46.17 ;
   RECT 23.18 46.17 508.44 47.88 ;
   RECT 23.18 47.88 508.44 49.59 ;
   RECT 23.18 49.59 508.44 51.3 ;
   RECT 23.18 51.3 508.44 53.01 ;
   RECT 23.18 53.01 508.44 54.72 ;
   RECT 23.18 54.72 508.44 56.43 ;
   RECT 23.18 56.43 508.44 58.14 ;
   RECT 23.18 58.14 508.44 59.85 ;
   RECT 23.18 59.85 508.44 61.56 ;
   RECT 23.18 61.56 508.44 63.27 ;
   RECT 23.18 63.27 508.44 64.98 ;
   RECT 23.18 64.98 508.44 66.69 ;
   RECT 23.18 66.69 508.44 68.4 ;
   RECT 23.18 68.4 508.44 70.11 ;
   RECT 23.18 70.11 508.44 71.82 ;
   RECT 23.18 71.82 508.44 73.53 ;
   RECT 23.18 73.53 508.44 75.24 ;
   RECT 23.18 75.24 508.44 76.95 ;
   RECT 23.18 76.95 508.44 78.66 ;
   RECT 23.18 78.66 508.44 80.37 ;
   RECT 23.18 80.37 508.44 82.08 ;
   RECT 23.18 82.08 508.44 83.79 ;
   RECT 23.18 83.79 508.44 85.5 ;
   RECT 23.18 85.5 508.44 87.21 ;
   RECT 23.18 87.21 508.44 88.92 ;
   RECT 23.18 88.92 508.44 90.63 ;
   RECT 23.18 90.63 508.44 92.34 ;
   RECT 23.18 92.34 508.44 94.05 ;
   RECT 23.18 94.05 508.44 95.76 ;
   RECT 23.18 95.76 508.44 97.47 ;
   RECT 23.18 97.47 508.44 99.18 ;
   RECT 23.18 99.18 508.44 100.89 ;
   RECT 23.18 100.89 508.44 102.6 ;
   RECT 23.18 102.6 508.44 104.31 ;
   RECT 23.18 104.31 508.44 106.02 ;
   RECT 23.18 106.02 508.44 107.73 ;
   RECT 23.18 107.73 508.44 109.44 ;
   RECT 23.18 109.44 508.44 111.15 ;
   RECT 23.18 111.15 508.44 112.86 ;
   RECT 23.18 112.86 508.44 114.57 ;
   RECT 23.18 114.57 508.44 116.28 ;
   RECT 23.18 116.28 508.44 117.99 ;
   RECT 23.18 117.99 508.44 119.7 ;
   RECT 23.18 119.7 508.44 121.41 ;
   RECT 23.18 121.41 508.44 123.12 ;
   RECT 23.18 123.12 508.44 124.83 ;
   RECT 23.18 124.83 508.44 126.54 ;
   RECT 23.18 126.54 508.44 128.25 ;
   RECT 23.18 128.25 508.44 129.96 ;
   RECT 23.18 129.96 508.44 131.67 ;
   RECT 23.18 131.67 508.44 133.38 ;
   RECT 23.18 133.38 508.44 135.09 ;
   RECT 23.18 135.09 508.44 136.8 ;
   RECT 23.18 136.8 508.44 138.51 ;
   RECT 23.18 138.51 508.44 140.22 ;
   RECT 23.18 140.22 508.44 141.93 ;
   RECT 23.18 141.93 508.44 143.64 ;
   RECT 23.18 143.64 508.44 145.35 ;
   RECT 23.18 145.35 508.44 147.06 ;
   RECT 23.18 147.06 508.44 148.77 ;
   RECT 23.18 148.77 508.44 150.48 ;
   RECT 0.0 150.48 508.44 152.19 ;
   RECT 0.0 152.19 508.44 153.9 ;
   RECT 0.0 153.9 508.44 155.61 ;
   RECT 0.0 155.61 508.44 157.32 ;
   RECT 0.0 157.32 508.44 159.03 ;
   RECT 0.0 159.03 508.44 160.74 ;
   RECT 0.0 160.74 508.44 162.45 ;
   RECT 0.0 162.45 508.44 164.16 ;
   RECT 0.0 164.16 508.44 165.87 ;
   RECT 0.0 165.87 508.44 167.58 ;
   RECT 0.0 167.58 508.44 169.29 ;
   RECT 0.0 169.29 508.44 171.0 ;
   RECT 0.0 171.0 508.44 172.71 ;
   RECT 0.0 172.71 508.44 174.42 ;
   RECT 0.0 174.42 508.44 176.13 ;
   RECT 0.0 176.13 508.44 177.84 ;
   RECT 0.0 177.84 508.44 179.55 ;
   RECT 23.18 179.55 508.44 181.26 ;
   RECT 23.18 181.26 508.44 182.97 ;
   RECT 23.18 182.97 508.44 184.68 ;
   RECT 23.18 184.68 508.44 186.39 ;
   RECT 23.18 186.39 508.44 188.1 ;
   RECT 23.18 188.1 508.44 189.81 ;
   RECT 23.18 189.81 508.44 191.52 ;
   RECT 23.18 191.52 508.44 193.23 ;
   RECT 23.18 193.23 508.44 194.94 ;
   RECT 23.18 194.94 508.44 196.65 ;
   RECT 23.18 196.65 508.44 198.36 ;
   RECT 23.18 198.36 508.44 200.07 ;
   RECT 23.18 200.07 508.44 201.78 ;
   RECT 23.18 201.78 508.44 203.49 ;
   RECT 23.18 203.49 508.44 205.2 ;
   RECT 23.18 205.2 508.44 206.91 ;
   RECT 23.18 206.91 508.44 208.62 ;
   RECT 23.18 208.62 508.44 210.33 ;
   RECT 23.18 210.33 508.44 212.04 ;
   RECT 23.18 212.04 508.44 213.75 ;
   RECT 23.18 213.75 508.44 215.46 ;
   RECT 23.18 215.46 508.44 217.17 ;
   RECT 23.18 217.17 508.44 218.88 ;
   RECT 23.18 218.88 508.44 220.59 ;
   RECT 23.18 220.59 508.44 222.3 ;
   RECT 23.18 222.3 508.44 224.01 ;
   RECT 23.18 224.01 508.44 225.72 ;
   RECT 23.18 225.72 508.44 227.43 ;
   RECT 23.18 227.43 508.44 229.14 ;
   RECT 23.18 229.14 508.44 230.85 ;
   RECT 23.18 230.85 508.44 232.56 ;
   RECT 23.18 232.56 508.44 234.27 ;
   RECT 23.18 234.27 508.44 235.98 ;
   RECT 23.18 235.98 508.44 237.69 ;
   RECT 23.18 237.69 508.44 239.4 ;
   RECT 23.18 239.4 508.44 241.11 ;
   RECT 23.18 241.11 508.44 242.82 ;
   RECT 23.18 242.82 508.44 244.53 ;
   RECT 23.18 244.53 508.44 246.24 ;
   RECT 23.18 246.24 508.44 247.95 ;
   RECT 23.18 247.95 508.44 249.66 ;
   RECT 23.18 249.66 508.44 251.37 ;
   RECT 23.18 251.37 508.44 253.08 ;
   RECT 23.18 253.08 508.44 254.79 ;
   RECT 23.18 254.79 508.44 256.5 ;
   RECT 23.18 256.5 508.44 258.21 ;
   RECT 23.18 258.21 508.44 259.92 ;
   RECT 23.18 259.92 508.44 261.63 ;
   RECT 23.18 261.63 508.44 263.34 ;
   RECT 23.18 263.34 508.44 265.05 ;
   RECT 23.18 265.05 508.44 266.76 ;
   RECT 23.18 266.76 508.44 268.47 ;
   RECT 23.18 268.47 508.44 270.18 ;
   RECT 23.18 270.18 508.44 271.89 ;
   RECT 23.18 271.89 508.44 273.6 ;
   RECT 23.18 273.6 508.44 275.31 ;
   RECT 23.18 275.31 508.44 277.02 ;
   RECT 23.18 277.02 508.44 278.73 ;
   RECT 23.18 278.73 508.44 280.44 ;
   RECT 23.18 280.44 508.44 282.15 ;
   RECT 23.18 282.15 508.44 283.86 ;
   RECT 23.18 283.86 508.44 285.57 ;
   RECT 23.18 285.57 508.44 287.28 ;
   RECT 23.18 287.28 508.44 288.99 ;
   RECT 23.18 288.99 508.44 290.7 ;
   RECT 23.18 290.7 508.44 292.41 ;
   RECT 23.18 292.41 508.44 294.12 ;
   RECT 23.18 294.12 508.44 295.83 ;
   RECT 23.18 295.83 508.44 297.54 ;
   RECT 23.18 297.54 508.44 299.25 ;
   RECT 23.18 299.25 508.44 300.96 ;
   RECT 23.18 300.96 508.44 302.67 ;
   RECT 23.18 302.67 508.44 304.38 ;
   RECT 23.18 304.38 508.44 306.09 ;
   RECT 23.18 306.09 508.44 307.8 ;
   RECT 23.18 307.8 508.44 309.51 ;
   RECT 23.18 309.51 508.44 311.22 ;
   RECT 23.18 311.22 508.44 312.93 ;
   RECT 23.18 312.93 508.44 314.64 ;
   RECT 23.18 314.64 508.44 316.35 ;
   RECT 23.18 316.35 508.44 318.06 ;
   RECT 23.18 318.06 508.44 319.77 ;
   RECT 23.18 319.77 508.44 321.48 ;
   RECT 23.18 321.48 508.44 323.19 ;
   RECT 23.18 323.19 508.44 324.9 ;
   RECT 23.18 324.9 508.44 326.61 ;
   RECT 23.18 326.61 508.44 328.32 ;
   RECT 23.18 328.32 508.44 330.03 ;
   RECT 23.18 330.03 508.44 331.74 ;
   RECT 23.18 331.74 508.44 333.45 ;
   RECT 23.18 333.45 508.44 335.16 ;
   RECT 23.18 335.16 508.44 336.87 ;
  LAYER metal3 ;
   RECT 23.18 0.0 508.44 1.71 ;
   RECT 23.18 1.71 508.44 3.42 ;
   RECT 23.18 3.42 508.44 5.13 ;
   RECT 23.18 5.13 508.44 6.84 ;
   RECT 23.18 6.84 508.44 8.55 ;
   RECT 23.18 8.55 508.44 10.26 ;
   RECT 23.18 10.26 508.44 11.97 ;
   RECT 23.18 11.97 508.44 13.68 ;
   RECT 23.18 13.68 508.44 15.39 ;
   RECT 23.18 15.39 508.44 17.1 ;
   RECT 23.18 17.1 508.44 18.81 ;
   RECT 23.18 18.81 508.44 20.52 ;
   RECT 23.18 20.52 508.44 22.23 ;
   RECT 23.18 22.23 508.44 23.94 ;
   RECT 23.18 23.94 508.44 25.65 ;
   RECT 23.18 25.65 508.44 27.36 ;
   RECT 23.18 27.36 508.44 29.07 ;
   RECT 23.18 29.07 508.44 30.78 ;
   RECT 23.18 30.78 508.44 32.49 ;
   RECT 23.18 32.49 508.44 34.2 ;
   RECT 23.18 34.2 508.44 35.91 ;
   RECT 23.18 35.91 508.44 37.62 ;
   RECT 23.18 37.62 508.44 39.33 ;
   RECT 23.18 39.33 508.44 41.04 ;
   RECT 23.18 41.04 508.44 42.75 ;
   RECT 23.18 42.75 508.44 44.46 ;
   RECT 23.18 44.46 508.44 46.17 ;
   RECT 23.18 46.17 508.44 47.88 ;
   RECT 23.18 47.88 508.44 49.59 ;
   RECT 23.18 49.59 508.44 51.3 ;
   RECT 23.18 51.3 508.44 53.01 ;
   RECT 23.18 53.01 508.44 54.72 ;
   RECT 23.18 54.72 508.44 56.43 ;
   RECT 23.18 56.43 508.44 58.14 ;
   RECT 23.18 58.14 508.44 59.85 ;
   RECT 23.18 59.85 508.44 61.56 ;
   RECT 23.18 61.56 508.44 63.27 ;
   RECT 23.18 63.27 508.44 64.98 ;
   RECT 23.18 64.98 508.44 66.69 ;
   RECT 23.18 66.69 508.44 68.4 ;
   RECT 23.18 68.4 508.44 70.11 ;
   RECT 23.18 70.11 508.44 71.82 ;
   RECT 23.18 71.82 508.44 73.53 ;
   RECT 23.18 73.53 508.44 75.24 ;
   RECT 23.18 75.24 508.44 76.95 ;
   RECT 23.18 76.95 508.44 78.66 ;
   RECT 23.18 78.66 508.44 80.37 ;
   RECT 23.18 80.37 508.44 82.08 ;
   RECT 23.18 82.08 508.44 83.79 ;
   RECT 23.18 83.79 508.44 85.5 ;
   RECT 23.18 85.5 508.44 87.21 ;
   RECT 23.18 87.21 508.44 88.92 ;
   RECT 23.18 88.92 508.44 90.63 ;
   RECT 23.18 90.63 508.44 92.34 ;
   RECT 23.18 92.34 508.44 94.05 ;
   RECT 23.18 94.05 508.44 95.76 ;
   RECT 23.18 95.76 508.44 97.47 ;
   RECT 23.18 97.47 508.44 99.18 ;
   RECT 23.18 99.18 508.44 100.89 ;
   RECT 23.18 100.89 508.44 102.6 ;
   RECT 23.18 102.6 508.44 104.31 ;
   RECT 23.18 104.31 508.44 106.02 ;
   RECT 23.18 106.02 508.44 107.73 ;
   RECT 23.18 107.73 508.44 109.44 ;
   RECT 23.18 109.44 508.44 111.15 ;
   RECT 23.18 111.15 508.44 112.86 ;
   RECT 23.18 112.86 508.44 114.57 ;
   RECT 23.18 114.57 508.44 116.28 ;
   RECT 23.18 116.28 508.44 117.99 ;
   RECT 23.18 117.99 508.44 119.7 ;
   RECT 23.18 119.7 508.44 121.41 ;
   RECT 23.18 121.41 508.44 123.12 ;
   RECT 23.18 123.12 508.44 124.83 ;
   RECT 23.18 124.83 508.44 126.54 ;
   RECT 23.18 126.54 508.44 128.25 ;
   RECT 23.18 128.25 508.44 129.96 ;
   RECT 23.18 129.96 508.44 131.67 ;
   RECT 23.18 131.67 508.44 133.38 ;
   RECT 23.18 133.38 508.44 135.09 ;
   RECT 23.18 135.09 508.44 136.8 ;
   RECT 23.18 136.8 508.44 138.51 ;
   RECT 23.18 138.51 508.44 140.22 ;
   RECT 23.18 140.22 508.44 141.93 ;
   RECT 23.18 141.93 508.44 143.64 ;
   RECT 23.18 143.64 508.44 145.35 ;
   RECT 23.18 145.35 508.44 147.06 ;
   RECT 23.18 147.06 508.44 148.77 ;
   RECT 23.18 148.77 508.44 150.48 ;
   RECT 0.0 150.48 508.44 152.19 ;
   RECT 0.0 152.19 508.44 153.9 ;
   RECT 0.0 153.9 508.44 155.61 ;
   RECT 0.0 155.61 508.44 157.32 ;
   RECT 0.0 157.32 508.44 159.03 ;
   RECT 0.0 159.03 508.44 160.74 ;
   RECT 0.0 160.74 508.44 162.45 ;
   RECT 0.0 162.45 508.44 164.16 ;
   RECT 0.0 164.16 508.44 165.87 ;
   RECT 0.0 165.87 508.44 167.58 ;
   RECT 0.0 167.58 508.44 169.29 ;
   RECT 0.0 169.29 508.44 171.0 ;
   RECT 0.0 171.0 508.44 172.71 ;
   RECT 0.0 172.71 508.44 174.42 ;
   RECT 0.0 174.42 508.44 176.13 ;
   RECT 0.0 176.13 508.44 177.84 ;
   RECT 0.0 177.84 508.44 179.55 ;
   RECT 23.18 179.55 508.44 181.26 ;
   RECT 23.18 181.26 508.44 182.97 ;
   RECT 23.18 182.97 508.44 184.68 ;
   RECT 23.18 184.68 508.44 186.39 ;
   RECT 23.18 186.39 508.44 188.1 ;
   RECT 23.18 188.1 508.44 189.81 ;
   RECT 23.18 189.81 508.44 191.52 ;
   RECT 23.18 191.52 508.44 193.23 ;
   RECT 23.18 193.23 508.44 194.94 ;
   RECT 23.18 194.94 508.44 196.65 ;
   RECT 23.18 196.65 508.44 198.36 ;
   RECT 23.18 198.36 508.44 200.07 ;
   RECT 23.18 200.07 508.44 201.78 ;
   RECT 23.18 201.78 508.44 203.49 ;
   RECT 23.18 203.49 508.44 205.2 ;
   RECT 23.18 205.2 508.44 206.91 ;
   RECT 23.18 206.91 508.44 208.62 ;
   RECT 23.18 208.62 508.44 210.33 ;
   RECT 23.18 210.33 508.44 212.04 ;
   RECT 23.18 212.04 508.44 213.75 ;
   RECT 23.18 213.75 508.44 215.46 ;
   RECT 23.18 215.46 508.44 217.17 ;
   RECT 23.18 217.17 508.44 218.88 ;
   RECT 23.18 218.88 508.44 220.59 ;
   RECT 23.18 220.59 508.44 222.3 ;
   RECT 23.18 222.3 508.44 224.01 ;
   RECT 23.18 224.01 508.44 225.72 ;
   RECT 23.18 225.72 508.44 227.43 ;
   RECT 23.18 227.43 508.44 229.14 ;
   RECT 23.18 229.14 508.44 230.85 ;
   RECT 23.18 230.85 508.44 232.56 ;
   RECT 23.18 232.56 508.44 234.27 ;
   RECT 23.18 234.27 508.44 235.98 ;
   RECT 23.18 235.98 508.44 237.69 ;
   RECT 23.18 237.69 508.44 239.4 ;
   RECT 23.18 239.4 508.44 241.11 ;
   RECT 23.18 241.11 508.44 242.82 ;
   RECT 23.18 242.82 508.44 244.53 ;
   RECT 23.18 244.53 508.44 246.24 ;
   RECT 23.18 246.24 508.44 247.95 ;
   RECT 23.18 247.95 508.44 249.66 ;
   RECT 23.18 249.66 508.44 251.37 ;
   RECT 23.18 251.37 508.44 253.08 ;
   RECT 23.18 253.08 508.44 254.79 ;
   RECT 23.18 254.79 508.44 256.5 ;
   RECT 23.18 256.5 508.44 258.21 ;
   RECT 23.18 258.21 508.44 259.92 ;
   RECT 23.18 259.92 508.44 261.63 ;
   RECT 23.18 261.63 508.44 263.34 ;
   RECT 23.18 263.34 508.44 265.05 ;
   RECT 23.18 265.05 508.44 266.76 ;
   RECT 23.18 266.76 508.44 268.47 ;
   RECT 23.18 268.47 508.44 270.18 ;
   RECT 23.18 270.18 508.44 271.89 ;
   RECT 23.18 271.89 508.44 273.6 ;
   RECT 23.18 273.6 508.44 275.31 ;
   RECT 23.18 275.31 508.44 277.02 ;
   RECT 23.18 277.02 508.44 278.73 ;
   RECT 23.18 278.73 508.44 280.44 ;
   RECT 23.18 280.44 508.44 282.15 ;
   RECT 23.18 282.15 508.44 283.86 ;
   RECT 23.18 283.86 508.44 285.57 ;
   RECT 23.18 285.57 508.44 287.28 ;
   RECT 23.18 287.28 508.44 288.99 ;
   RECT 23.18 288.99 508.44 290.7 ;
   RECT 23.18 290.7 508.44 292.41 ;
   RECT 23.18 292.41 508.44 294.12 ;
   RECT 23.18 294.12 508.44 295.83 ;
   RECT 23.18 295.83 508.44 297.54 ;
   RECT 23.18 297.54 508.44 299.25 ;
   RECT 23.18 299.25 508.44 300.96 ;
   RECT 23.18 300.96 508.44 302.67 ;
   RECT 23.18 302.67 508.44 304.38 ;
   RECT 23.18 304.38 508.44 306.09 ;
   RECT 23.18 306.09 508.44 307.8 ;
   RECT 23.18 307.8 508.44 309.51 ;
   RECT 23.18 309.51 508.44 311.22 ;
   RECT 23.18 311.22 508.44 312.93 ;
   RECT 23.18 312.93 508.44 314.64 ;
   RECT 23.18 314.64 508.44 316.35 ;
   RECT 23.18 316.35 508.44 318.06 ;
   RECT 23.18 318.06 508.44 319.77 ;
   RECT 23.18 319.77 508.44 321.48 ;
   RECT 23.18 321.48 508.44 323.19 ;
   RECT 23.18 323.19 508.44 324.9 ;
   RECT 23.18 324.9 508.44 326.61 ;
   RECT 23.18 326.61 508.44 328.32 ;
   RECT 23.18 328.32 508.44 330.03 ;
   RECT 23.18 330.03 508.44 331.74 ;
   RECT 23.18 331.74 508.44 333.45 ;
   RECT 23.18 333.45 508.44 335.16 ;
   RECT 23.18 335.16 508.44 336.87 ;
  LAYER via3 ;
   RECT 23.18 0.0 508.44 1.71 ;
   RECT 23.18 1.71 508.44 3.42 ;
   RECT 23.18 3.42 508.44 5.13 ;
   RECT 23.18 5.13 508.44 6.84 ;
   RECT 23.18 6.84 508.44 8.55 ;
   RECT 23.18 8.55 508.44 10.26 ;
   RECT 23.18 10.26 508.44 11.97 ;
   RECT 23.18 11.97 508.44 13.68 ;
   RECT 23.18 13.68 508.44 15.39 ;
   RECT 23.18 15.39 508.44 17.1 ;
   RECT 23.18 17.1 508.44 18.81 ;
   RECT 23.18 18.81 508.44 20.52 ;
   RECT 23.18 20.52 508.44 22.23 ;
   RECT 23.18 22.23 508.44 23.94 ;
   RECT 23.18 23.94 508.44 25.65 ;
   RECT 23.18 25.65 508.44 27.36 ;
   RECT 23.18 27.36 508.44 29.07 ;
   RECT 23.18 29.07 508.44 30.78 ;
   RECT 23.18 30.78 508.44 32.49 ;
   RECT 23.18 32.49 508.44 34.2 ;
   RECT 23.18 34.2 508.44 35.91 ;
   RECT 23.18 35.91 508.44 37.62 ;
   RECT 23.18 37.62 508.44 39.33 ;
   RECT 23.18 39.33 508.44 41.04 ;
   RECT 23.18 41.04 508.44 42.75 ;
   RECT 23.18 42.75 508.44 44.46 ;
   RECT 23.18 44.46 508.44 46.17 ;
   RECT 23.18 46.17 508.44 47.88 ;
   RECT 23.18 47.88 508.44 49.59 ;
   RECT 23.18 49.59 508.44 51.3 ;
   RECT 23.18 51.3 508.44 53.01 ;
   RECT 23.18 53.01 508.44 54.72 ;
   RECT 23.18 54.72 508.44 56.43 ;
   RECT 23.18 56.43 508.44 58.14 ;
   RECT 23.18 58.14 508.44 59.85 ;
   RECT 23.18 59.85 508.44 61.56 ;
   RECT 23.18 61.56 508.44 63.27 ;
   RECT 23.18 63.27 508.44 64.98 ;
   RECT 23.18 64.98 508.44 66.69 ;
   RECT 23.18 66.69 508.44 68.4 ;
   RECT 23.18 68.4 508.44 70.11 ;
   RECT 23.18 70.11 508.44 71.82 ;
   RECT 23.18 71.82 508.44 73.53 ;
   RECT 23.18 73.53 508.44 75.24 ;
   RECT 23.18 75.24 508.44 76.95 ;
   RECT 23.18 76.95 508.44 78.66 ;
   RECT 23.18 78.66 508.44 80.37 ;
   RECT 23.18 80.37 508.44 82.08 ;
   RECT 23.18 82.08 508.44 83.79 ;
   RECT 23.18 83.79 508.44 85.5 ;
   RECT 23.18 85.5 508.44 87.21 ;
   RECT 23.18 87.21 508.44 88.92 ;
   RECT 23.18 88.92 508.44 90.63 ;
   RECT 23.18 90.63 508.44 92.34 ;
   RECT 23.18 92.34 508.44 94.05 ;
   RECT 23.18 94.05 508.44 95.76 ;
   RECT 23.18 95.76 508.44 97.47 ;
   RECT 23.18 97.47 508.44 99.18 ;
   RECT 23.18 99.18 508.44 100.89 ;
   RECT 23.18 100.89 508.44 102.6 ;
   RECT 23.18 102.6 508.44 104.31 ;
   RECT 23.18 104.31 508.44 106.02 ;
   RECT 23.18 106.02 508.44 107.73 ;
   RECT 23.18 107.73 508.44 109.44 ;
   RECT 23.18 109.44 508.44 111.15 ;
   RECT 23.18 111.15 508.44 112.86 ;
   RECT 23.18 112.86 508.44 114.57 ;
   RECT 23.18 114.57 508.44 116.28 ;
   RECT 23.18 116.28 508.44 117.99 ;
   RECT 23.18 117.99 508.44 119.7 ;
   RECT 23.18 119.7 508.44 121.41 ;
   RECT 23.18 121.41 508.44 123.12 ;
   RECT 23.18 123.12 508.44 124.83 ;
   RECT 23.18 124.83 508.44 126.54 ;
   RECT 23.18 126.54 508.44 128.25 ;
   RECT 23.18 128.25 508.44 129.96 ;
   RECT 23.18 129.96 508.44 131.67 ;
   RECT 23.18 131.67 508.44 133.38 ;
   RECT 23.18 133.38 508.44 135.09 ;
   RECT 23.18 135.09 508.44 136.8 ;
   RECT 23.18 136.8 508.44 138.51 ;
   RECT 23.18 138.51 508.44 140.22 ;
   RECT 23.18 140.22 508.44 141.93 ;
   RECT 23.18 141.93 508.44 143.64 ;
   RECT 23.18 143.64 508.44 145.35 ;
   RECT 23.18 145.35 508.44 147.06 ;
   RECT 23.18 147.06 508.44 148.77 ;
   RECT 23.18 148.77 508.44 150.48 ;
   RECT 0.0 150.48 508.44 152.19 ;
   RECT 0.0 152.19 508.44 153.9 ;
   RECT 0.0 153.9 508.44 155.61 ;
   RECT 0.0 155.61 508.44 157.32 ;
   RECT 0.0 157.32 508.44 159.03 ;
   RECT 0.0 159.03 508.44 160.74 ;
   RECT 0.0 160.74 508.44 162.45 ;
   RECT 0.0 162.45 508.44 164.16 ;
   RECT 0.0 164.16 508.44 165.87 ;
   RECT 0.0 165.87 508.44 167.58 ;
   RECT 0.0 167.58 508.44 169.29 ;
   RECT 0.0 169.29 508.44 171.0 ;
   RECT 0.0 171.0 508.44 172.71 ;
   RECT 0.0 172.71 508.44 174.42 ;
   RECT 0.0 174.42 508.44 176.13 ;
   RECT 0.0 176.13 508.44 177.84 ;
   RECT 0.0 177.84 508.44 179.55 ;
   RECT 23.18 179.55 508.44 181.26 ;
   RECT 23.18 181.26 508.44 182.97 ;
   RECT 23.18 182.97 508.44 184.68 ;
   RECT 23.18 184.68 508.44 186.39 ;
   RECT 23.18 186.39 508.44 188.1 ;
   RECT 23.18 188.1 508.44 189.81 ;
   RECT 23.18 189.81 508.44 191.52 ;
   RECT 23.18 191.52 508.44 193.23 ;
   RECT 23.18 193.23 508.44 194.94 ;
   RECT 23.18 194.94 508.44 196.65 ;
   RECT 23.18 196.65 508.44 198.36 ;
   RECT 23.18 198.36 508.44 200.07 ;
   RECT 23.18 200.07 508.44 201.78 ;
   RECT 23.18 201.78 508.44 203.49 ;
   RECT 23.18 203.49 508.44 205.2 ;
   RECT 23.18 205.2 508.44 206.91 ;
   RECT 23.18 206.91 508.44 208.62 ;
   RECT 23.18 208.62 508.44 210.33 ;
   RECT 23.18 210.33 508.44 212.04 ;
   RECT 23.18 212.04 508.44 213.75 ;
   RECT 23.18 213.75 508.44 215.46 ;
   RECT 23.18 215.46 508.44 217.17 ;
   RECT 23.18 217.17 508.44 218.88 ;
   RECT 23.18 218.88 508.44 220.59 ;
   RECT 23.18 220.59 508.44 222.3 ;
   RECT 23.18 222.3 508.44 224.01 ;
   RECT 23.18 224.01 508.44 225.72 ;
   RECT 23.18 225.72 508.44 227.43 ;
   RECT 23.18 227.43 508.44 229.14 ;
   RECT 23.18 229.14 508.44 230.85 ;
   RECT 23.18 230.85 508.44 232.56 ;
   RECT 23.18 232.56 508.44 234.27 ;
   RECT 23.18 234.27 508.44 235.98 ;
   RECT 23.18 235.98 508.44 237.69 ;
   RECT 23.18 237.69 508.44 239.4 ;
   RECT 23.18 239.4 508.44 241.11 ;
   RECT 23.18 241.11 508.44 242.82 ;
   RECT 23.18 242.82 508.44 244.53 ;
   RECT 23.18 244.53 508.44 246.24 ;
   RECT 23.18 246.24 508.44 247.95 ;
   RECT 23.18 247.95 508.44 249.66 ;
   RECT 23.18 249.66 508.44 251.37 ;
   RECT 23.18 251.37 508.44 253.08 ;
   RECT 23.18 253.08 508.44 254.79 ;
   RECT 23.18 254.79 508.44 256.5 ;
   RECT 23.18 256.5 508.44 258.21 ;
   RECT 23.18 258.21 508.44 259.92 ;
   RECT 23.18 259.92 508.44 261.63 ;
   RECT 23.18 261.63 508.44 263.34 ;
   RECT 23.18 263.34 508.44 265.05 ;
   RECT 23.18 265.05 508.44 266.76 ;
   RECT 23.18 266.76 508.44 268.47 ;
   RECT 23.18 268.47 508.44 270.18 ;
   RECT 23.18 270.18 508.44 271.89 ;
   RECT 23.18 271.89 508.44 273.6 ;
   RECT 23.18 273.6 508.44 275.31 ;
   RECT 23.18 275.31 508.44 277.02 ;
   RECT 23.18 277.02 508.44 278.73 ;
   RECT 23.18 278.73 508.44 280.44 ;
   RECT 23.18 280.44 508.44 282.15 ;
   RECT 23.18 282.15 508.44 283.86 ;
   RECT 23.18 283.86 508.44 285.57 ;
   RECT 23.18 285.57 508.44 287.28 ;
   RECT 23.18 287.28 508.44 288.99 ;
   RECT 23.18 288.99 508.44 290.7 ;
   RECT 23.18 290.7 508.44 292.41 ;
   RECT 23.18 292.41 508.44 294.12 ;
   RECT 23.18 294.12 508.44 295.83 ;
   RECT 23.18 295.83 508.44 297.54 ;
   RECT 23.18 297.54 508.44 299.25 ;
   RECT 23.18 299.25 508.44 300.96 ;
   RECT 23.18 300.96 508.44 302.67 ;
   RECT 23.18 302.67 508.44 304.38 ;
   RECT 23.18 304.38 508.44 306.09 ;
   RECT 23.18 306.09 508.44 307.8 ;
   RECT 23.18 307.8 508.44 309.51 ;
   RECT 23.18 309.51 508.44 311.22 ;
   RECT 23.18 311.22 508.44 312.93 ;
   RECT 23.18 312.93 508.44 314.64 ;
   RECT 23.18 314.64 508.44 316.35 ;
   RECT 23.18 316.35 508.44 318.06 ;
   RECT 23.18 318.06 508.44 319.77 ;
   RECT 23.18 319.77 508.44 321.48 ;
   RECT 23.18 321.48 508.44 323.19 ;
   RECT 23.18 323.19 508.44 324.9 ;
   RECT 23.18 324.9 508.44 326.61 ;
   RECT 23.18 326.61 508.44 328.32 ;
   RECT 23.18 328.32 508.44 330.03 ;
   RECT 23.18 330.03 508.44 331.74 ;
   RECT 23.18 331.74 508.44 333.45 ;
   RECT 23.18 333.45 508.44 335.16 ;
   RECT 23.18 335.16 508.44 336.87 ;
  LAYER metal4 ;
   RECT 23.18 0.0 508.44 1.71 ;
   RECT 23.18 1.71 508.44 3.42 ;
   RECT 23.18 3.42 508.44 5.13 ;
   RECT 23.18 5.13 508.44 6.84 ;
   RECT 23.18 6.84 508.44 8.55 ;
   RECT 23.18 8.55 508.44 10.26 ;
   RECT 23.18 10.26 508.44 11.97 ;
   RECT 23.18 11.97 508.44 13.68 ;
   RECT 23.18 13.68 508.44 15.39 ;
   RECT 23.18 15.39 508.44 17.1 ;
   RECT 23.18 17.1 508.44 18.81 ;
   RECT 23.18 18.81 508.44 20.52 ;
   RECT 23.18 20.52 508.44 22.23 ;
   RECT 23.18 22.23 508.44 23.94 ;
   RECT 23.18 23.94 508.44 25.65 ;
   RECT 23.18 25.65 508.44 27.36 ;
   RECT 23.18 27.36 508.44 29.07 ;
   RECT 23.18 29.07 508.44 30.78 ;
   RECT 23.18 30.78 508.44 32.49 ;
   RECT 23.18 32.49 508.44 34.2 ;
   RECT 23.18 34.2 508.44 35.91 ;
   RECT 23.18 35.91 508.44 37.62 ;
   RECT 23.18 37.62 508.44 39.33 ;
   RECT 23.18 39.33 508.44 41.04 ;
   RECT 23.18 41.04 508.44 42.75 ;
   RECT 23.18 42.75 508.44 44.46 ;
   RECT 23.18 44.46 508.44 46.17 ;
   RECT 23.18 46.17 508.44 47.88 ;
   RECT 23.18 47.88 508.44 49.59 ;
   RECT 23.18 49.59 508.44 51.3 ;
   RECT 23.18 51.3 508.44 53.01 ;
   RECT 23.18 53.01 508.44 54.72 ;
   RECT 23.18 54.72 508.44 56.43 ;
   RECT 23.18 56.43 508.44 58.14 ;
   RECT 23.18 58.14 508.44 59.85 ;
   RECT 23.18 59.85 508.44 61.56 ;
   RECT 23.18 61.56 508.44 63.27 ;
   RECT 23.18 63.27 508.44 64.98 ;
   RECT 23.18 64.98 508.44 66.69 ;
   RECT 23.18 66.69 508.44 68.4 ;
   RECT 23.18 68.4 508.44 70.11 ;
   RECT 23.18 70.11 508.44 71.82 ;
   RECT 23.18 71.82 508.44 73.53 ;
   RECT 23.18 73.53 508.44 75.24 ;
   RECT 23.18 75.24 508.44 76.95 ;
   RECT 23.18 76.95 508.44 78.66 ;
   RECT 23.18 78.66 508.44 80.37 ;
   RECT 23.18 80.37 508.44 82.08 ;
   RECT 23.18 82.08 508.44 83.79 ;
   RECT 23.18 83.79 508.44 85.5 ;
   RECT 23.18 85.5 508.44 87.21 ;
   RECT 23.18 87.21 508.44 88.92 ;
   RECT 23.18 88.92 508.44 90.63 ;
   RECT 23.18 90.63 508.44 92.34 ;
   RECT 23.18 92.34 508.44 94.05 ;
   RECT 23.18 94.05 508.44 95.76 ;
   RECT 23.18 95.76 508.44 97.47 ;
   RECT 23.18 97.47 508.44 99.18 ;
   RECT 23.18 99.18 508.44 100.89 ;
   RECT 23.18 100.89 508.44 102.6 ;
   RECT 23.18 102.6 508.44 104.31 ;
   RECT 23.18 104.31 508.44 106.02 ;
   RECT 23.18 106.02 508.44 107.73 ;
   RECT 23.18 107.73 508.44 109.44 ;
   RECT 23.18 109.44 508.44 111.15 ;
   RECT 23.18 111.15 508.44 112.86 ;
   RECT 23.18 112.86 508.44 114.57 ;
   RECT 23.18 114.57 508.44 116.28 ;
   RECT 23.18 116.28 508.44 117.99 ;
   RECT 23.18 117.99 508.44 119.7 ;
   RECT 23.18 119.7 508.44 121.41 ;
   RECT 23.18 121.41 508.44 123.12 ;
   RECT 23.18 123.12 508.44 124.83 ;
   RECT 23.18 124.83 508.44 126.54 ;
   RECT 23.18 126.54 508.44 128.25 ;
   RECT 23.18 128.25 508.44 129.96 ;
   RECT 23.18 129.96 508.44 131.67 ;
   RECT 23.18 131.67 508.44 133.38 ;
   RECT 23.18 133.38 508.44 135.09 ;
   RECT 23.18 135.09 508.44 136.8 ;
   RECT 23.18 136.8 508.44 138.51 ;
   RECT 23.18 138.51 508.44 140.22 ;
   RECT 23.18 140.22 508.44 141.93 ;
   RECT 23.18 141.93 508.44 143.64 ;
   RECT 23.18 143.64 508.44 145.35 ;
   RECT 23.18 145.35 508.44 147.06 ;
   RECT 23.18 147.06 508.44 148.77 ;
   RECT 23.18 148.77 508.44 150.48 ;
   RECT 0.0 150.48 508.44 152.19 ;
   RECT 0.0 152.19 508.44 153.9 ;
   RECT 0.0 153.9 508.44 155.61 ;
   RECT 0.0 155.61 508.44 157.32 ;
   RECT 0.0 157.32 508.44 159.03 ;
   RECT 0.0 159.03 508.44 160.74 ;
   RECT 0.0 160.74 508.44 162.45 ;
   RECT 0.0 162.45 508.44 164.16 ;
   RECT 0.0 164.16 508.44 165.87 ;
   RECT 0.0 165.87 508.44 167.58 ;
   RECT 0.0 167.58 508.44 169.29 ;
   RECT 0.0 169.29 508.44 171.0 ;
   RECT 0.0 171.0 508.44 172.71 ;
   RECT 0.0 172.71 508.44 174.42 ;
   RECT 0.0 174.42 508.44 176.13 ;
   RECT 0.0 176.13 508.44 177.84 ;
   RECT 0.0 177.84 508.44 179.55 ;
   RECT 23.18 179.55 508.44 181.26 ;
   RECT 23.18 181.26 508.44 182.97 ;
   RECT 23.18 182.97 508.44 184.68 ;
   RECT 23.18 184.68 508.44 186.39 ;
   RECT 23.18 186.39 508.44 188.1 ;
   RECT 23.18 188.1 508.44 189.81 ;
   RECT 23.18 189.81 508.44 191.52 ;
   RECT 23.18 191.52 508.44 193.23 ;
   RECT 23.18 193.23 508.44 194.94 ;
   RECT 23.18 194.94 508.44 196.65 ;
   RECT 23.18 196.65 508.44 198.36 ;
   RECT 23.18 198.36 508.44 200.07 ;
   RECT 23.18 200.07 508.44 201.78 ;
   RECT 23.18 201.78 508.44 203.49 ;
   RECT 23.18 203.49 508.44 205.2 ;
   RECT 23.18 205.2 508.44 206.91 ;
   RECT 23.18 206.91 508.44 208.62 ;
   RECT 23.18 208.62 508.44 210.33 ;
   RECT 23.18 210.33 508.44 212.04 ;
   RECT 23.18 212.04 508.44 213.75 ;
   RECT 23.18 213.75 508.44 215.46 ;
   RECT 23.18 215.46 508.44 217.17 ;
   RECT 23.18 217.17 508.44 218.88 ;
   RECT 23.18 218.88 508.44 220.59 ;
   RECT 23.18 220.59 508.44 222.3 ;
   RECT 23.18 222.3 508.44 224.01 ;
   RECT 23.18 224.01 508.44 225.72 ;
   RECT 23.18 225.72 508.44 227.43 ;
   RECT 23.18 227.43 508.44 229.14 ;
   RECT 23.18 229.14 508.44 230.85 ;
   RECT 23.18 230.85 508.44 232.56 ;
   RECT 23.18 232.56 508.44 234.27 ;
   RECT 23.18 234.27 508.44 235.98 ;
   RECT 23.18 235.98 508.44 237.69 ;
   RECT 23.18 237.69 508.44 239.4 ;
   RECT 23.18 239.4 508.44 241.11 ;
   RECT 23.18 241.11 508.44 242.82 ;
   RECT 23.18 242.82 508.44 244.53 ;
   RECT 23.18 244.53 508.44 246.24 ;
   RECT 23.18 246.24 508.44 247.95 ;
   RECT 23.18 247.95 508.44 249.66 ;
   RECT 23.18 249.66 508.44 251.37 ;
   RECT 23.18 251.37 508.44 253.08 ;
   RECT 23.18 253.08 508.44 254.79 ;
   RECT 23.18 254.79 508.44 256.5 ;
   RECT 23.18 256.5 508.44 258.21 ;
   RECT 23.18 258.21 508.44 259.92 ;
   RECT 23.18 259.92 508.44 261.63 ;
   RECT 23.18 261.63 508.44 263.34 ;
   RECT 23.18 263.34 508.44 265.05 ;
   RECT 23.18 265.05 508.44 266.76 ;
   RECT 23.18 266.76 508.44 268.47 ;
   RECT 23.18 268.47 508.44 270.18 ;
   RECT 23.18 270.18 508.44 271.89 ;
   RECT 23.18 271.89 508.44 273.6 ;
   RECT 23.18 273.6 508.44 275.31 ;
   RECT 23.18 275.31 508.44 277.02 ;
   RECT 23.18 277.02 508.44 278.73 ;
   RECT 23.18 278.73 508.44 280.44 ;
   RECT 23.18 280.44 508.44 282.15 ;
   RECT 23.18 282.15 508.44 283.86 ;
   RECT 23.18 283.86 508.44 285.57 ;
   RECT 23.18 285.57 508.44 287.28 ;
   RECT 23.18 287.28 508.44 288.99 ;
   RECT 23.18 288.99 508.44 290.7 ;
   RECT 23.18 290.7 508.44 292.41 ;
   RECT 23.18 292.41 508.44 294.12 ;
   RECT 23.18 294.12 508.44 295.83 ;
   RECT 23.18 295.83 508.44 297.54 ;
   RECT 23.18 297.54 508.44 299.25 ;
   RECT 23.18 299.25 508.44 300.96 ;
   RECT 23.18 300.96 508.44 302.67 ;
   RECT 23.18 302.67 508.44 304.38 ;
   RECT 23.18 304.38 508.44 306.09 ;
   RECT 23.18 306.09 508.44 307.8 ;
   RECT 23.18 307.8 508.44 309.51 ;
   RECT 23.18 309.51 508.44 311.22 ;
   RECT 23.18 311.22 508.44 312.93 ;
   RECT 23.18 312.93 508.44 314.64 ;
   RECT 23.18 314.64 508.44 316.35 ;
   RECT 23.18 316.35 508.44 318.06 ;
   RECT 23.18 318.06 508.44 319.77 ;
   RECT 23.18 319.77 508.44 321.48 ;
   RECT 23.18 321.48 508.44 323.19 ;
   RECT 23.18 323.19 508.44 324.9 ;
   RECT 23.18 324.9 508.44 326.61 ;
   RECT 23.18 326.61 508.44 328.32 ;
   RECT 23.18 328.32 508.44 330.03 ;
   RECT 23.18 330.03 508.44 331.74 ;
   RECT 23.18 331.74 508.44 333.45 ;
   RECT 23.18 333.45 508.44 335.16 ;
   RECT 23.18 335.16 508.44 336.87 ;
 END
END block_1338x1773_192

MACRO block_546x684_100
 CLASS BLOCK ;
 FOREIGN block_546x684_100 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 207.48 BY 129.96 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.135 126.825 117.705 127.395 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 4.275 3.325 4.845 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 20.995 3.325 21.565 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 20.235 3.325 20.805 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 18.715 3.325 19.285 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 62.035 3.325 62.605 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 58.995 3.325 59.565 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 58.235 3.325 58.805 ;
  END
 END o7
 PIN o8
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 110.675 126.825 111.245 127.395 ;
  END
 END o8
 PIN o9
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 107.255 126.825 107.825 127.395 ;
  END
 END o9
 PIN o10
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 119.795 126.825 120.365 127.395 ;
  END
 END o10
 PIN o11
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 18.335 204.345 18.905 ;
  END
 END o11
 PIN o12
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 19.855 204.345 20.425 ;
  END
 END o12
 PIN o13
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 20.615 204.345 21.185 ;
  END
 END o13
 PIN o14
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 21.375 204.345 21.945 ;
  END
 END o14
 PIN o15
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 22.135 204.345 22.705 ;
  END
 END o15
 PIN o16
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 22.895 204.345 23.465 ;
  END
 END o16
 PIN o17
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 24.415 204.345 24.985 ;
  END
 END o17
 PIN o18
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 25.175 204.345 25.745 ;
  END
 END o18
 PIN o19
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 25.935 204.345 26.505 ;
  END
 END o19
 PIN o20
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 26.695 204.345 27.265 ;
  END
 END o20
 PIN o21
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 27.455 204.345 28.025 ;
  END
 END o21
 PIN o22
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 28.975 204.345 29.545 ;
  END
 END o22
 PIN o23
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 29.735 204.345 30.305 ;
  END
 END o23
 PIN o24
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 30.495 204.345 31.065 ;
  END
 END o24
 PIN o25
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 31.255 204.345 31.825 ;
  END
 END o25
 PIN o26
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 48.735 204.345 49.305 ;
  END
 END o26
 PIN o27
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 33.535 204.345 34.105 ;
  END
 END o27
 PIN o28
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.325 80.56 174.895 81.13 ;
  END
 END o28
 PIN o29
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 35.055 204.345 35.625 ;
  END
 END o29
 PIN o30
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 35.815 204.345 36.385 ;
  END
 END o30
 PIN o31
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 36.575 204.345 37.145 ;
  END
 END o31
 PIN o32
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 38.095 204.345 38.665 ;
  END
 END o32
 PIN o33
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 38.855 204.345 39.425 ;
  END
 END o33
 PIN o34
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 39.615 204.345 40.185 ;
  END
 END o34
 PIN o35
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 40.375 204.345 40.945 ;
  END
 END o35
 PIN o36
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 41.135 204.345 41.705 ;
  END
 END o36
 PIN o37
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 42.655 204.345 43.225 ;
  END
 END o37
 PIN o38
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 43.415 204.345 43.985 ;
  END
 END o38
 PIN o39
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 44.175 204.345 44.745 ;
  END
 END o39
 PIN o40
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 44.935 204.345 45.505 ;
  END
 END o40
 PIN o41
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 45.695 204.345 46.265 ;
  END
 END o41
 PIN o42
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 47.215 204.345 47.785 ;
  END
 END o42
 PIN o43
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 47.975 204.345 48.545 ;
  END
 END o43
 PIN o44
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 49.495 204.345 50.065 ;
  END
 END o44
 PIN o45
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 50.255 204.345 50.825 ;
  END
 END o45
 PIN o46
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 51.775 204.345 52.345 ;
  END
 END o46
 PIN o47
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 52.535 204.345 53.105 ;
  END
 END o47
 PIN o48
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 53.295 204.345 53.865 ;
  END
 END o48
 PIN o49
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 54.055 204.345 54.625 ;
  END
 END o49
 PIN o50
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 54.815 204.345 55.385 ;
  END
 END o50
 PIN o51
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 95.095 126.825 95.665 127.395 ;
  END
 END o51
 PIN o52
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 101.555 126.825 102.125 127.395 ;
  END
 END o52
 PIN o53
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 104.215 126.825 104.785 127.395 ;
  END
 END o53
 PIN o54
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 114.095 126.825 114.665 127.395 ;
  END
 END o54
 PIN o55
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 132.715 126.825 133.285 127.395 ;
  END
 END o55
 PIN o56
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 153.995 126.825 154.565 127.395 ;
  END
 END o56
 PIN o57
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 172.995 126.825 173.565 127.395 ;
  END
 END o57
 PIN o58
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 176.035 126.825 176.605 127.395 ;
  END
 END o58
 PIN o59
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 179.455 126.825 180.025 127.395 ;
  END
 END o59
 PIN o60
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 181.735 126.825 182.305 127.395 ;
  END
 END o60
 PIN o61
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 185.155 126.825 185.725 127.395 ;
  END
 END o61
 PIN o62
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 188.575 126.825 189.145 127.395 ;
  END
 END o62
 PIN o63
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 200.735 126.825 201.305 127.395 ;
  END
 END o63
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 82.935 126.825 83.505 127.395 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 70.395 126.825 70.965 127.395 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 85.975 126.825 86.545 127.395 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 41.895 126.825 42.465 127.395 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 44.935 126.825 45.505 127.395 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 48.355 126.825 48.925 127.395 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 51.775 126.825 52.345 127.395 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 54.815 126.825 55.385 127.395 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 57.475 126.825 58.045 127.395 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 60.515 126.825 61.085 127.395 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 63.935 126.825 64.505 127.395 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 88.635 126.825 89.205 127.395 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 73.055 126.825 73.625 127.395 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 91.675 126.825 92.245 127.395 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 98.515 126.825 99.085 127.395 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 126.825 130.245 127.395 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 150.955 126.825 151.525 127.395 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 197.315 126.825 197.885 127.395 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 77.995 3.325 78.565 ;
  END
 END i18
 PIN i19
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 76.475 3.325 77.045 ;
  END
 END i19
 PIN i20
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 75.715 3.325 76.285 ;
  END
 END i20
 PIN i21
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 79.515 3.325 80.085 ;
  END
 END i21
 PIN i22
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 56.335 204.345 56.905 ;
  END
 END i22
 PIN i23
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 57.095 204.345 57.665 ;
  END
 END i23
 PIN i24
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 57.855 204.345 58.425 ;
  END
 END i24
 PIN i25
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 58.615 204.345 59.185 ;
  END
 END i25
 PIN i26
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 59.375 204.345 59.945 ;
  END
 END i26
 PIN i27
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 60.895 204.345 61.465 ;
  END
 END i27
 PIN i28
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 63.175 204.345 63.745 ;
  END
 END i28
 PIN i29
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 63.935 204.345 64.505 ;
  END
 END i29
 PIN i30
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 65.455 204.345 66.025 ;
  END
 END i30
 PIN i31
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 66.215 204.345 66.785 ;
  END
 END i31
 PIN i32
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 66.975 204.345 67.545 ;
  END
 END i32
 PIN i33
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.775 67.735 204.345 68.305 ;
  END
 END i33
 PIN i34
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 74.955 3.325 75.525 ;
  END
 END i34
 PIN i35
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 77.235 3.325 77.805 ;
  END
 END i35
 OBS
  LAYER metal1 ;
   RECT 0 0 207.48 129.96 ;
  LAYER via1 ;
   RECT 0 0 207.48 129.96 ;
  LAYER metal2 ;
   RECT 0 0 207.48 129.96 ;
  LAYER via2 ;
   RECT 0 0 207.48 129.96 ;
  LAYER metal3 ;
   RECT 0 0 207.48 129.96 ;
  LAYER via3 ;
   RECT 0 0 207.48 129.96 ;
  LAYER metal4 ;
   RECT 0 0 207.48 129.96 ;
 END
END block_546x684_100

MACRO block_737x1152_453
 CLASS BLOCK ;
 FOREIGN block_737x1152_453 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 280.06 BY 218.88 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 93.955 0.855 94.525 1.425 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 96.995 0.855 97.565 1.425 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 100.035 0.855 100.605 1.425 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 103.075 0.855 103.645 1.425 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 106.115 0.855 106.685 1.425 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 109.155 0.855 109.725 1.425 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 112.195 0.855 112.765 1.425 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 115.235 0.855 115.805 1.425 ;
  END
 END o7
 PIN o8
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 32.395 0.855 32.965 1.425 ;
  END
 END o8
 PIN o9
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 35.435 0.855 36.005 1.425 ;
  END
 END o9
 PIN o10
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 38.475 0.855 39.045 1.425 ;
  END
 END o10
 PIN o11
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 41.515 0.855 42.085 1.425 ;
  END
 END o11
 PIN o12
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 44.555 0.855 45.125 1.425 ;
  END
 END o12
 PIN o13
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 47.595 0.855 48.165 1.425 ;
  END
 END o13
 PIN o14
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 50.635 0.855 51.205 1.425 ;
  END
 END o14
 PIN o15
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 53.675 0.855 54.245 1.425 ;
  END
 END o15
 PIN o16
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 119.795 0.855 120.365 1.425 ;
  END
 END o16
 PIN o17
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 122.835 0.855 123.405 1.425 ;
  END
 END o17
 PIN o18
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 0.855 126.445 1.425 ;
  END
 END o18
 PIN o19
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 128.915 0.855 129.485 1.425 ;
  END
 END o19
 PIN o20
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 131.955 0.855 132.525 1.425 ;
  END
 END o20
 PIN o21
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 134.995 0.855 135.565 1.425 ;
  END
 END o21
 PIN o22
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 138.035 0.855 138.605 1.425 ;
  END
 END o22
 PIN o23
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 141.075 0.855 141.645 1.425 ;
  END
 END o23
 PIN o24
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 6.555 0.855 7.125 1.425 ;
  END
 END o24
 PIN o25
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.595 0.855 10.165 1.425 ;
  END
 END o25
 PIN o26
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 12.635 0.855 13.205 1.425 ;
  END
 END o26
 PIN o27
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 15.675 0.855 16.245 1.425 ;
  END
 END o27
 PIN o28
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 18.715 0.855 19.285 1.425 ;
  END
 END o28
 PIN o29
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 21.755 0.855 22.325 1.425 ;
  END
 END o29
 PIN o30
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 24.795 0.855 25.365 1.425 ;
  END
 END o30
 PIN o31
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 0.855 28.405 1.425 ;
  END
 END o31
 PIN o32
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 61.655 251.465 62.225 ;
  END
 END o32
 PIN o33
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 66.025 251.465 66.595 ;
  END
 END o33
 PIN o34
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 64.695 251.465 65.265 ;
  END
 END o34
 PIN o35
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 20.995 251.465 21.565 ;
  END
 END o35
 PIN o36
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 39.805 251.465 40.375 ;
  END
 END o36
 PIN o37
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 34.105 251.465 34.675 ;
  END
 END o37
 PIN o38
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 25.365 251.465 25.935 ;
  END
 END o38
 PIN o39
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 38.475 251.465 39.045 ;
  END
 END o39
 PIN o40
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 31.065 251.465 31.635 ;
  END
 END o40
 PIN o41
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 42.845 251.465 43.415 ;
  END
 END o41
 PIN o42
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 44.175 251.465 44.745 ;
  END
 END o42
 PIN o43
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 35.435 251.465 36.005 ;
  END
 END o43
 PIN o44
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 29.735 251.465 30.305 ;
  END
 END o44
 PIN o45
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 22.325 251.465 22.895 ;
  END
 END o45
 PIN o46
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 26.695 251.465 27.265 ;
  END
 END o46
 PIN o47
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 60.325 251.465 60.895 ;
  END
 END o47
 PIN o48
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 55.955 251.465 56.525 ;
  END
 END o48
 PIN o49
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 51.585 251.465 52.155 ;
  END
 END o49
 PIN o50
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 47.215 251.465 47.785 ;
  END
 END o50
 PIN o51
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 108.395 251.465 108.965 ;
  END
 END o51
 PIN o52
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 77.805 251.465 78.375 ;
  END
 END o52
 PIN o53
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 112.765 251.465 113.335 ;
  END
 END o53
 PIN o54
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 131.575 251.465 132.145 ;
  END
 END o54
 PIN o55
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 92.245 251.465 92.815 ;
  END
 END o55
 PIN o56
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 121.505 251.465 122.075 ;
  END
 END o56
 PIN o57
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 127.205 251.465 127.775 ;
  END
 END o57
 PIN o58
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 109.725 251.465 110.295 ;
  END
 END o58
 PIN o59
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 79.135 251.465 79.705 ;
  END
 END o59
 PIN o60
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 130.245 251.465 130.815 ;
  END
 END o60
 PIN o61
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 125.875 251.465 126.445 ;
  END
 END o61
 PIN o62
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 122.835 251.465 123.405 ;
  END
 END o62
 PIN o63
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 117.135 251.465 117.705 ;
  END
 END o63
 PIN o64
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 114.095 251.465 114.665 ;
  END
 END o64
 PIN o65
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 73.435 251.465 74.005 ;
  END
 END o65
 PIN o66
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 70.395 251.465 70.965 ;
  END
 END o66
 PIN o67
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 74.765 251.465 75.335 ;
  END
 END o67
 PIN o68
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 118.465 251.465 119.035 ;
  END
 END o68
 PIN o69
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 69.065 251.465 69.635 ;
  END
 END o69
 PIN o70
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 83.505 251.465 84.075 ;
  END
 END o70
 PIN o71
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 86.545 251.465 87.115 ;
  END
 END o71
 PIN o72
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 95.285 251.465 95.855 ;
  END
 END o72
 PIN o73
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 87.875 251.465 88.445 ;
  END
 END o73
 PIN o74
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 82.175 251.465 82.745 ;
  END
 END o74
 PIN o75
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 90.915 251.465 91.485 ;
  END
 END o75
 PIN o76
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 105.355 251.465 105.925 ;
  END
 END o76
 PIN o77
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 104.025 251.465 104.595 ;
  END
 END o77
 PIN o78
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 100.985 251.465 101.555 ;
  END
 END o78
 PIN o79
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 168.435 251.465 169.005 ;
  END
 END o79
 PIN o80
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 99.655 251.465 100.225 ;
  END
 END o80
 PIN o81
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 96.615 251.465 97.185 ;
  END
 END o81
 PIN o82
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 170.715 251.465 171.285 ;
  END
 END o82
 PIN o83
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 48.545 251.465 49.115 ;
  END
 END o83
 PIN o84
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 52.915 251.465 53.485 ;
  END
 END o84
 PIN o85
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.895 57.285 251.465 57.855 ;
  END
 END o85
 PIN o86
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 139.935 0.855 140.505 1.425 ;
  END
 END o86
 PIN o87
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 130.815 0.855 131.385 1.425 ;
  END
 END o87
 PIN o88
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 104.975 0.855 105.545 1.425 ;
  END
 END o88
 PIN o89
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 114.095 0.855 114.665 1.425 ;
  END
 END o89
 PIN o90
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 101.935 0.855 102.505 1.425 ;
  END
 END o90
 PIN o91
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 133.855 0.855 134.425 1.425 ;
  END
 END o91
 PIN o92
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 111.055 0.855 111.625 1.425 ;
  END
 END o92
 PIN o93
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 95.855 0.855 96.425 1.425 ;
  END
 END o93
 PIN o94
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.135 0.855 117.705 1.425 ;
  END
 END o94
 PIN o95
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 124.735 0.855 125.305 1.425 ;
  END
 END o95
 PIN o96
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 127.775 0.855 128.345 1.425 ;
  END
 END o96
 PIN o97
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 98.895 0.855 99.465 1.425 ;
  END
 END o97
 PIN o98
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 121.695 0.855 122.265 1.425 ;
  END
 END o98
 PIN o99
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 52.535 0.855 53.105 1.425 ;
  END
 END o99
 PIN o100
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 40.375 0.855 40.945 1.425 ;
  END
 END o100
 PIN o101
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 17.575 0.855 18.145 1.425 ;
  END
 END o101
 PIN o102
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 49.495 0.855 50.065 1.425 ;
  END
 END o102
 PIN o103
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 37.335 0.855 37.905 1.425 ;
  END
 END o103
 PIN o104
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 0.855 27.265 1.425 ;
  END
 END o104
 PIN o105
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 14.535 0.855 15.105 1.425 ;
  END
 END o105
 PIN o106
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.295 0.855 34.865 1.425 ;
  END
 END o106
 PIN o107
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 46.455 0.855 47.025 1.425 ;
  END
 END o107
 PIN o108
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 8.455 0.855 9.025 1.425 ;
  END
 END o108
 PIN o109
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 43.415 0.855 43.985 1.425 ;
  END
 END o109
 PIN o110
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 11.495 0.855 12.065 1.425 ;
  END
 END o110
 PIN o111
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 20.615 0.855 21.185 1.425 ;
  END
 END o111
 PIN o112
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 29.735 0.855 30.305 1.425 ;
  END
 END o112
 PIN o113
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 136.895 0.855 137.465 1.425 ;
  END
 END o113
 PIN o114
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 23.655 0.855 24.225 1.425 ;
  END
 END o114
 PIN o115
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.575 0.855 56.145 1.425 ;
  END
 END o115
 PIN o116
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 142.975 0.855 143.545 1.425 ;
  END
 END o116
 PIN o117
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 108.015 0.855 108.585 1.425 ;
  END
 END o117
 PIN o118
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 74.195 0.855 74.765 1.425 ;
  END
 END o118
 PIN o119
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 207.575 216.885 208.145 217.455 ;
  END
 END o119
 PIN o120
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 250.135 0.855 250.705 1.425 ;
  END
 END o120
 PIN o121
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 170.145 277.305 170.715 ;
  END
 END o121
 PIN o122
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 169.385 277.305 169.955 ;
  END
 END o122
 PIN o123
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 113.905 277.305 114.475 ;
  END
 END o123
 PIN o124
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 113.145 277.305 113.715 ;
  END
 END o124
 PIN o125
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 109.535 277.305 110.105 ;
  END
 END o125
 PIN o126
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 108.775 277.305 109.345 ;
  END
 END o126
 PIN o127
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 105.165 277.305 105.735 ;
  END
 END o127
 PIN o128
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 104.405 277.305 104.975 ;
  END
 END o128
 PIN o129
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 100.795 277.305 101.365 ;
  END
 END o129
 PIN o130
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 100.035 277.305 100.605 ;
  END
 END o130
 PIN o131
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 96.425 277.305 96.995 ;
  END
 END o131
 PIN o132
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 95.665 277.305 96.235 ;
  END
 END o132
 PIN o133
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 131.385 277.305 131.955 ;
  END
 END o133
 PIN o134
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 92.055 277.305 92.625 ;
  END
 END o134
 PIN o135
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 91.295 277.305 91.865 ;
  END
 END o135
 PIN o136
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 87.685 277.305 88.255 ;
  END
 END o136
 PIN o137
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 86.925 277.305 87.495 ;
  END
 END o137
 PIN o138
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 83.315 277.305 83.885 ;
  END
 END o138
 PIN o139
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 82.555 277.305 83.125 ;
  END
 END o139
 PIN o140
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 78.945 277.305 79.515 ;
  END
 END o140
 PIN o141
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 78.185 277.305 78.755 ;
  END
 END o141
 PIN o142
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 74.575 277.305 75.145 ;
  END
 END o142
 PIN o143
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 73.815 277.305 74.385 ;
  END
 END o143
 PIN o144
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 130.625 277.305 131.195 ;
  END
 END o144
 PIN o145
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 70.205 277.305 70.775 ;
  END
 END o145
 PIN o146
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 69.445 277.305 70.015 ;
  END
 END o146
 PIN o147
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 65.835 277.305 66.405 ;
  END
 END o147
 PIN o148
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 65.075 277.305 65.645 ;
  END
 END o148
 PIN o149
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 61.465 277.305 62.035 ;
  END
 END o149
 PIN o150
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 60.705 277.305 61.275 ;
  END
 END o150
 PIN o151
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 57.095 277.305 57.665 ;
  END
 END o151
 PIN o152
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 56.335 277.305 56.905 ;
  END
 END o152
 PIN o153
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 52.725 277.305 53.295 ;
  END
 END o153
 PIN o154
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 51.965 277.305 52.535 ;
  END
 END o154
 PIN o155
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 127.015 277.305 127.585 ;
  END
 END o155
 PIN o156
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 48.355 277.305 48.925 ;
  END
 END o156
 PIN o157
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 47.595 277.305 48.165 ;
  END
 END o157
 PIN o158
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 43.985 277.305 44.555 ;
  END
 END o158
 PIN o159
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 43.225 277.305 43.795 ;
  END
 END o159
 PIN o160
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 39.615 277.305 40.185 ;
  END
 END o160
 PIN o161
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 38.855 277.305 39.425 ;
  END
 END o161
 PIN o162
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 35.245 277.305 35.815 ;
  END
 END o162
 PIN o163
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 34.485 277.305 35.055 ;
  END
 END o163
 PIN o164
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 30.875 277.305 31.445 ;
  END
 END o164
 PIN o165
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 30.115 277.305 30.685 ;
  END
 END o165
 PIN o166
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 126.255 277.305 126.825 ;
  END
 END o166
 PIN o167
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 26.505 277.305 27.075 ;
  END
 END o167
 PIN o168
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 25.745 277.305 26.315 ;
  END
 END o168
 PIN o169
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 22.135 277.305 22.705 ;
  END
 END o169
 PIN o170
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 21.375 277.305 21.945 ;
  END
 END o170
 PIN o171
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 122.645 277.305 123.215 ;
  END
 END o171
 PIN o172
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 121.885 277.305 122.455 ;
  END
 END o172
 PIN o173
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 118.275 277.305 118.845 ;
  END
 END o173
 PIN o174
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 117.515 277.305 118.085 ;
  END
 END o174
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 235.315 216.885 235.885 217.455 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 224.675 216.885 225.245 217.455 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 223.915 216.885 224.485 217.455 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 237.215 216.885 237.785 217.455 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 223.155 216.885 223.725 217.455 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 236.075 216.885 236.645 217.455 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 123.215 269.705 123.785 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 121.125 269.705 121.695 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 118.845 269.705 119.415 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 116.755 269.705 117.325 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 114.475 269.705 115.045 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 112.385 269.705 112.955 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 129.865 269.705 130.435 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 127.585 269.705 128.155 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 125.495 269.705 126.065 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 170.525 269.705 171.095 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 168.435 269.705 169.005 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 131.955 269.705 132.525 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 75.145 269.705 75.715 ;
  END
 END i18
 PIN i19
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 73.055 269.705 73.625 ;
  END
 END i19
 PIN i20
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 70.775 269.705 71.345 ;
  END
 END i20
 PIN i21
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 68.685 269.705 69.255 ;
  END
 END i21
 PIN i22
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 66.405 269.705 66.975 ;
  END
 END i22
 PIN i23
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 64.315 269.705 64.885 ;
  END
 END i23
 PIN i24
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 83.885 269.705 84.455 ;
  END
 END i24
 PIN i25
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 81.795 269.705 82.365 ;
  END
 END i25
 PIN i26
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 79.515 269.705 80.085 ;
  END
 END i26
 PIN i27
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 77.425 269.705 77.995 ;
  END
 END i27
 PIN i28
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 38.095 269.705 38.665 ;
  END
 END i28
 PIN i29
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 35.815 269.705 36.385 ;
  END
 END i29
 PIN i30
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 33.725 269.705 34.295 ;
  END
 END i30
 PIN i31
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 31.445 269.705 32.015 ;
  END
 END i31
 PIN i32
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 29.355 269.705 29.925 ;
  END
 END i32
 PIN i33
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 27.075 269.705 27.645 ;
  END
 END i33
 PIN i34
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 24.985 269.705 25.555 ;
  END
 END i34
 PIN i35
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 22.705 269.705 23.275 ;
  END
 END i35
 PIN i36
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 20.615 269.705 21.185 ;
  END
 END i36
 PIN i37
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 62.035 269.705 62.605 ;
  END
 END i37
 PIN i38
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 59.945 269.705 60.515 ;
  END
 END i38
 PIN i39
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 57.665 269.705 58.235 ;
  END
 END i39
 PIN i40
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 55.575 269.705 56.145 ;
  END
 END i40
 PIN i41
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 53.295 269.705 53.865 ;
  END
 END i41
 PIN i42
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 51.205 269.705 51.775 ;
  END
 END i42
 PIN i43
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 48.925 269.705 49.495 ;
  END
 END i43
 PIN i44
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 46.835 269.705 47.405 ;
  END
 END i44
 PIN i45
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 44.555 269.705 45.125 ;
  END
 END i45
 PIN i46
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 42.465 269.705 43.035 ;
  END
 END i46
 PIN i47
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 40.185 269.705 40.755 ;
  END
 END i47
 PIN i48
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 110.105 269.705 110.675 ;
  END
 END i48
 PIN i49
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 92.625 269.705 93.195 ;
  END
 END i49
 PIN i50
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 90.535 269.705 91.105 ;
  END
 END i50
 PIN i51
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 88.255 269.705 88.825 ;
  END
 END i51
 PIN i52
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 86.165 269.705 86.735 ;
  END
 END i52
 PIN i53
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 108.015 269.705 108.585 ;
  END
 END i53
 PIN i54
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 105.735 269.705 106.305 ;
  END
 END i54
 PIN i55
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 103.645 269.705 104.215 ;
  END
 END i55
 PIN i56
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 101.365 269.705 101.935 ;
  END
 END i56
 PIN i57
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 99.275 269.705 99.845 ;
  END
 END i57
 PIN i58
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 96.995 269.705 97.565 ;
  END
 END i58
 PIN i59
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.135 94.905 269.705 95.475 ;
  END
 END i59
 PIN i60
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 220.115 216.885 220.685 217.455 ;
  END
 END i60
 PIN i61
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.775 216.885 242.345 217.455 ;
  END
 END i61
 PIN i62
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 243.675 216.885 244.245 217.455 ;
  END
 END i62
 PIN i63
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 218.595 216.885 219.165 217.455 ;
  END
 END i63
 PIN i64
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 239.875 216.885 240.445 217.455 ;
  END
 END i64
 PIN i65
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 245.195 216.885 245.765 217.455 ;
  END
 END i65
 PIN i66
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 209.475 216.885 210.045 217.455 ;
  END
 END i66
 PIN i67
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 208.335 216.885 208.905 217.455 ;
  END
 END i67
 PIN i68
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.635 216.885 241.205 217.455 ;
  END
 END i68
 PIN i69
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 217.455 216.885 218.025 217.455 ;
  END
 END i69
 PIN i70
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 219.355 216.885 219.925 217.455 ;
  END
 END i70
 PIN i71
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 244.435 216.885 245.005 217.455 ;
  END
 END i71
 PIN i72
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 242.535 216.885 243.105 217.455 ;
  END
 END i72
 PIN i73
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 170.525 276.545 171.095 ;
  END
 END i73
 PIN i74
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 168.815 276.545 169.385 ;
  END
 END i74
 PIN i75
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 114.285 276.545 114.855 ;
  END
 END i75
 PIN i76
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 112.575 276.545 113.145 ;
  END
 END i76
 PIN i77
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 109.915 276.545 110.485 ;
  END
 END i77
 PIN i78
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 108.205 276.545 108.775 ;
  END
 END i78
 PIN i79
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 105.545 276.545 106.115 ;
  END
 END i79
 PIN i80
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 103.835 276.545 104.405 ;
  END
 END i80
 PIN i81
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 101.175 276.545 101.745 ;
  END
 END i81
 PIN i82
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 99.465 276.545 100.035 ;
  END
 END i82
 PIN i83
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 96.805 276.545 97.375 ;
  END
 END i83
 PIN i84
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 95.095 276.545 95.665 ;
  END
 END i84
 PIN i85
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 131.765 276.545 132.335 ;
  END
 END i85
 PIN i86
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 92.435 276.545 93.005 ;
  END
 END i86
 PIN i87
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 90.725 276.545 91.295 ;
  END
 END i87
 PIN i88
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 88.065 276.545 88.635 ;
  END
 END i88
 PIN i89
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 86.355 276.545 86.925 ;
  END
 END i89
 PIN i90
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 83.695 276.545 84.265 ;
  END
 END i90
 PIN i91
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 81.985 276.545 82.555 ;
  END
 END i91
 PIN i92
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 79.325 276.545 79.895 ;
  END
 END i92
 PIN i93
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 77.615 276.545 78.185 ;
  END
 END i93
 PIN i94
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 74.955 276.545 75.525 ;
  END
 END i94
 PIN i95
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 73.245 276.545 73.815 ;
  END
 END i95
 PIN i96
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 130.055 276.545 130.625 ;
  END
 END i96
 PIN i97
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 70.585 276.545 71.155 ;
  END
 END i97
 PIN i98
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 68.875 276.545 69.445 ;
  END
 END i98
 PIN i99
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 66.215 276.545 66.785 ;
  END
 END i99
 PIN i100
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 64.505 276.545 65.075 ;
  END
 END i100
 PIN i101
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 61.845 276.545 62.415 ;
  END
 END i101
 PIN i102
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 60.135 276.545 60.705 ;
  END
 END i102
 PIN i103
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 57.475 276.545 58.045 ;
  END
 END i103
 PIN i104
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 55.765 276.545 56.335 ;
  END
 END i104
 PIN i105
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 53.105 276.545 53.675 ;
  END
 END i105
 PIN i106
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 51.395 276.545 51.965 ;
  END
 END i106
 PIN i107
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 127.395 276.545 127.965 ;
  END
 END i107
 PIN i108
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 48.735 276.545 49.305 ;
  END
 END i108
 PIN i109
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 47.025 276.545 47.595 ;
  END
 END i109
 PIN i110
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 44.365 276.545 44.935 ;
  END
 END i110
 PIN i111
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 42.655 276.545 43.225 ;
  END
 END i111
 PIN i112
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 39.995 276.545 40.565 ;
  END
 END i112
 PIN i113
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 38.285 276.545 38.855 ;
  END
 END i113
 PIN i114
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 35.625 276.545 36.195 ;
  END
 END i114
 PIN i115
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 33.915 276.545 34.485 ;
  END
 END i115
 PIN i116
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 31.255 276.545 31.825 ;
  END
 END i116
 PIN i117
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 29.545 276.545 30.115 ;
  END
 END i117
 PIN i118
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 125.685 276.545 126.255 ;
  END
 END i118
 PIN i119
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 26.885 276.545 27.455 ;
  END
 END i119
 PIN i120
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 25.175 276.545 25.745 ;
  END
 END i120
 PIN i121
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 22.515 276.545 23.085 ;
  END
 END i121
 PIN i122
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 20.805 276.545 21.375 ;
  END
 END i122
 PIN i123
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 123.025 276.545 123.595 ;
  END
 END i123
 PIN i124
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 121.315 276.545 121.885 ;
  END
 END i124
 PIN i125
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 118.655 276.545 119.225 ;
  END
 END i125
 PIN i126
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 116.945 276.545 117.515 ;
  END
 END i126
 PIN i127
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 171.095 277.305 171.665 ;
  END
 END i127
 PIN i128
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 168.435 277.305 169.005 ;
  END
 END i128
 PIN i129
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 114.855 277.305 115.425 ;
  END
 END i129
 PIN i130
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 112.195 277.305 112.765 ;
  END
 END i130
 PIN i131
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 110.485 277.305 111.055 ;
  END
 END i131
 PIN i132
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 107.825 277.305 108.395 ;
  END
 END i132
 PIN i133
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 106.115 277.305 106.685 ;
  END
 END i133
 PIN i134
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 103.455 277.305 104.025 ;
  END
 END i134
 PIN i135
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 101.745 277.305 102.315 ;
  END
 END i135
 PIN i136
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 99.085 277.305 99.655 ;
  END
 END i136
 PIN i137
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 97.375 277.305 97.945 ;
  END
 END i137
 PIN i138
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 94.715 277.305 95.285 ;
  END
 END i138
 PIN i139
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 132.335 277.305 132.905 ;
  END
 END i139
 PIN i140
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 93.005 277.305 93.575 ;
  END
 END i140
 PIN i141
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 90.345 277.305 90.915 ;
  END
 END i141
 PIN i142
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 88.635 277.305 89.205 ;
  END
 END i142
 PIN i143
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 85.975 277.305 86.545 ;
  END
 END i143
 PIN i144
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 84.265 277.305 84.835 ;
  END
 END i144
 PIN i145
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 81.605 277.305 82.175 ;
  END
 END i145
 PIN i146
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 79.895 277.305 80.465 ;
  END
 END i146
 PIN i147
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 77.235 277.305 77.805 ;
  END
 END i147
 PIN i148
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 75.525 277.305 76.095 ;
  END
 END i148
 PIN i149
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 72.865 277.305 73.435 ;
  END
 END i149
 PIN i150
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 129.675 277.305 130.245 ;
  END
 END i150
 PIN i151
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 71.155 277.305 71.725 ;
  END
 END i151
 PIN i152
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 68.495 277.305 69.065 ;
  END
 END i152
 PIN i153
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 66.785 277.305 67.355 ;
  END
 END i153
 PIN i154
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 64.125 277.305 64.695 ;
  END
 END i154
 PIN i155
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 62.415 277.305 62.985 ;
  END
 END i155
 PIN i156
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 59.755 277.305 60.325 ;
  END
 END i156
 PIN i157
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 58.045 277.305 58.615 ;
  END
 END i157
 PIN i158
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 55.385 277.305 55.955 ;
  END
 END i158
 PIN i159
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 53.675 277.305 54.245 ;
  END
 END i159
 PIN i160
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 51.015 277.305 51.585 ;
  END
 END i160
 PIN i161
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 127.965 277.305 128.535 ;
  END
 END i161
 PIN i162
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 49.305 277.305 49.875 ;
  END
 END i162
 PIN i163
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 46.645 277.305 47.215 ;
  END
 END i163
 PIN i164
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 44.935 277.305 45.505 ;
  END
 END i164
 PIN i165
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 42.275 277.305 42.845 ;
  END
 END i165
 PIN i166
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 40.565 277.305 41.135 ;
  END
 END i166
 PIN i167
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 37.905 277.305 38.475 ;
  END
 END i167
 PIN i168
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 36.195 277.305 36.765 ;
  END
 END i168
 PIN i169
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 33.535 277.305 34.105 ;
  END
 END i169
 PIN i170
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 31.825 277.305 32.395 ;
  END
 END i170
 PIN i171
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 29.165 277.305 29.735 ;
  END
 END i171
 PIN i172
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 125.305 277.305 125.875 ;
  END
 END i172
 PIN i173
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 27.455 277.305 28.025 ;
  END
 END i173
 PIN i174
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 24.795 277.305 25.365 ;
  END
 END i174
 PIN i175
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 23.085 277.305 23.655 ;
  END
 END i175
 PIN i176
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 20.425 277.305 20.995 ;
  END
 END i176
 PIN i177
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 123.595 277.305 124.165 ;
  END
 END i177
 PIN i178
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 120.935 277.305 121.505 ;
  END
 END i178
 PIN i179
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 119.225 277.305 119.795 ;
  END
 END i179
 PIN i180
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 116.565 277.305 117.135 ;
  END
 END i180
 PIN i181
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 276.735 152.095 277.305 152.665 ;
  END
 END i181
 PIN i182
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 171.475 276.545 172.045 ;
  END
 END i182
 PIN i183
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 167.865 276.545 168.435 ;
  END
 END i183
 PIN i184
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 115.235 276.545 115.805 ;
  END
 END i184
 PIN i185
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 111.625 276.545 112.195 ;
  END
 END i185
 PIN i186
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 110.865 276.545 111.435 ;
  END
 END i186
 PIN i187
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 107.255 276.545 107.825 ;
  END
 END i187
 PIN i188
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 106.495 276.545 107.065 ;
  END
 END i188
 PIN i189
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 102.885 276.545 103.455 ;
  END
 END i189
 PIN i190
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 102.125 276.545 102.695 ;
  END
 END i190
 PIN i191
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 98.515 276.545 99.085 ;
  END
 END i191
 PIN i192
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 97.755 276.545 98.325 ;
  END
 END i192
 PIN i193
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 94.145 276.545 94.715 ;
  END
 END i193
 PIN i194
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 132.715 276.545 133.285 ;
  END
 END i194
 PIN i195
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 93.385 276.545 93.955 ;
  END
 END i195
 PIN i196
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 89.775 276.545 90.345 ;
  END
 END i196
 PIN i197
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 89.015 276.545 89.585 ;
  END
 END i197
 PIN i198
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 85.405 276.545 85.975 ;
  END
 END i198
 PIN i199
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 84.645 276.545 85.215 ;
  END
 END i199
 PIN i200
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 81.035 276.545 81.605 ;
  END
 END i200
 PIN i201
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 80.275 276.545 80.845 ;
  END
 END i201
 PIN i202
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 76.665 276.545 77.235 ;
  END
 END i202
 PIN i203
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 75.905 276.545 76.475 ;
  END
 END i203
 PIN i204
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 72.295 276.545 72.865 ;
  END
 END i204
 PIN i205
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 129.105 276.545 129.675 ;
  END
 END i205
 PIN i206
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 71.535 276.545 72.105 ;
  END
 END i206
 PIN i207
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 67.925 276.545 68.495 ;
  END
 END i207
 PIN i208
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 67.165 276.545 67.735 ;
  END
 END i208
 PIN i209
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 63.555 276.545 64.125 ;
  END
 END i209
 PIN i210
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 62.795 276.545 63.365 ;
  END
 END i210
 PIN i211
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 59.185 276.545 59.755 ;
  END
 END i211
 PIN i212
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 58.425 276.545 58.995 ;
  END
 END i212
 PIN i213
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 54.815 276.545 55.385 ;
  END
 END i213
 PIN i214
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 54.055 276.545 54.625 ;
  END
 END i214
 PIN i215
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 50.445 276.545 51.015 ;
  END
 END i215
 PIN i216
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 128.345 276.545 128.915 ;
  END
 END i216
 PIN i217
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 49.685 276.545 50.255 ;
  END
 END i217
 PIN i218
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 46.075 276.545 46.645 ;
  END
 END i218
 PIN i219
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 45.315 276.545 45.885 ;
  END
 END i219
 PIN i220
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 41.705 276.545 42.275 ;
  END
 END i220
 PIN i221
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 40.945 276.545 41.515 ;
  END
 END i221
 PIN i222
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 37.335 276.545 37.905 ;
  END
 END i222
 PIN i223
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 36.575 276.545 37.145 ;
  END
 END i223
 PIN i224
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 32.965 276.545 33.535 ;
  END
 END i224
 PIN i225
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 32.205 276.545 32.775 ;
  END
 END i225
 PIN i226
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 28.595 276.545 29.165 ;
  END
 END i226
 PIN i227
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 124.735 276.545 125.305 ;
  END
 END i227
 PIN i228
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 27.835 276.545 28.405 ;
  END
 END i228
 PIN i229
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 24.225 276.545 24.795 ;
  END
 END i229
 PIN i230
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 23.465 276.545 24.035 ;
  END
 END i230
 PIN i231
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 19.855 276.545 20.425 ;
  END
 END i231
 PIN i232
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 123.975 276.545 124.545 ;
  END
 END i232
 PIN i233
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 120.365 276.545 120.935 ;
  END
 END i233
 PIN i234
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 119.605 276.545 120.175 ;
  END
 END i234
 PIN i235
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 275.975 115.995 276.545 116.565 ;
  END
 END i235
 PIN i236
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 210.235 216.885 210.805 217.455 ;
  END
 END i236
 PIN i237
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 215.555 216.885 216.125 217.455 ;
  END
 END i237
 PIN i238
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 214.795 216.885 215.365 217.455 ;
  END
 END i238
 PIN i239
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 214.035 216.885 214.605 217.455 ;
  END
 END i239
 PIN i240
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 212.895 216.885 213.465 217.455 ;
  END
 END i240
 PIN i241
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 212.135 216.885 212.705 217.455 ;
  END
 END i241
 PIN i242
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 210.995 216.885 211.565 217.455 ;
  END
 END i242
 PIN i243
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 204.915 216.885 205.485 217.455 ;
  END
 END i243
 PIN i244
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 234.555 216.885 235.125 217.455 ;
  END
 END i244
 PIN i245
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 225.815 216.885 226.385 217.455 ;
  END
 END i245
 PIN i246
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 233.415 216.885 233.985 217.455 ;
  END
 END i246
 PIN i247
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 226.575 216.885 227.145 217.455 ;
  END
 END i247
 PIN i248
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 232.655 216.885 233.225 217.455 ;
  END
 END i248
 PIN i249
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 227.715 216.885 228.285 217.455 ;
  END
 END i249
 PIN i250
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 178.315 216.885 178.885 217.455 ;
  END
 END i250
 PIN i251
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.895 216.885 175.465 217.455 ;
  END
 END i251
 PIN i252
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 159.315 216.885 159.885 217.455 ;
  END
 END i252
 PIN i253
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.755 216.885 155.325 217.455 ;
  END
 END i253
 PIN i254
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 152.855 216.885 153.425 217.455 ;
  END
 END i254
 PIN i255
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 150.195 216.885 150.765 217.455 ;
  END
 END i255
 PIN i256
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 148.295 216.885 148.865 217.455 ;
  END
 END i256
 PIN i257
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 183.635 216.885 184.205 217.455 ;
  END
 END i257
 PIN i258
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 186.675 216.885 187.245 217.455 ;
  END
 END i258
 PIN i259
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 189.335 216.885 189.905 217.455 ;
  END
 END i259
 PIN i260
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 193.895 216.885 194.465 217.455 ;
  END
 END i260
 PIN i261
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 160.075 216.885 160.645 217.455 ;
  END
 END i261
 PIN i262
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 170.335 216.885 170.905 217.455 ;
  END
 END i262
 PIN i263
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 166.535 216.885 167.105 217.455 ;
  END
 END i263
 PIN i264
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 162.735 216.885 163.305 217.455 ;
  END
 END i264
 PIN i265
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 167.295 216.885 167.865 217.455 ;
  END
 END i265
 PIN i266
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 171.095 216.885 171.665 217.455 ;
  END
 END i266
 PIN i267
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.655 216.885 176.225 217.455 ;
  END
 END i267
 PIN i268
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 179.455 216.885 180.025 217.455 ;
  END
 END i268
 PIN i269
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 163.875 216.885 164.445 217.455 ;
  END
 END i269
 PIN i270
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 201.495 216.885 202.065 217.455 ;
  END
 END i270
 PIN i271
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 200.355 216.885 200.925 217.455 ;
  END
 END i271
 PIN i272
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 197.695 216.885 198.265 217.455 ;
  END
 END i272
 PIN i273
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 196.555 216.885 197.125 217.455 ;
  END
 END i273
 PIN i274
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 193.135 216.885 193.705 217.455 ;
  END
 END i274
 PIN i275
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 191.995 216.885 192.565 217.455 ;
  END
 END i275
 PIN i276
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 190.475 216.885 191.045 217.455 ;
  END
 END i276
 PIN i277
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 203.395 216.885 203.965 217.455 ;
  END
 END i277
 OBS
  LAYER metal1 ;
   RECT 0 0 280.06 218.88 ;
  LAYER via1 ;
   RECT 0 0 280.06 218.88 ;
  LAYER metal2 ;
   RECT 0 0 280.06 218.88 ;
  LAYER via2 ;
   RECT 0 0 280.06 218.88 ;
  LAYER metal3 ;
   RECT 0 0 280.06 218.88 ;
  LAYER via3 ;
   RECT 0 0 280.06 218.88 ;
  LAYER metal4 ;
   RECT 0 0 280.06 218.88 ;
 END
END block_737x1152_453

MACRO block_644x666_91
 CLASS BLOCK ;
 FOREIGN block_644x666_91 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 244.72 BY 126.54 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 33.535 241.585 34.105 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 33.915 240.825 34.485 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 34.295 241.585 34.865 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 34.675 240.825 35.245 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 35.055 241.585 35.625 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 35.435 240.825 36.005 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 35.815 241.585 36.385 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 36.195 240.825 36.765 ;
  END
 END o7
 PIN o8
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 36.575 241.585 37.145 ;
  END
 END o8
 PIN o9
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 36.955 240.825 37.525 ;
  END
 END o9
 PIN o10
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 38.095 241.585 38.665 ;
  END
 END o10
 PIN o11
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 38.475 240.825 39.045 ;
  END
 END o11
 PIN o12
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 38.855 241.585 39.425 ;
  END
 END o12
 PIN o13
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 39.235 240.825 39.805 ;
  END
 END o13
 PIN o14
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 39.615 241.585 40.185 ;
  END
 END o14
 PIN o15
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 39.995 240.825 40.565 ;
  END
 END o15
 PIN o16
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 40.375 241.585 40.945 ;
  END
 END o16
 PIN o17
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 40.755 240.825 41.325 ;
  END
 END o17
 PIN o18
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 41.135 241.585 41.705 ;
  END
 END o18
 PIN o19
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 43.415 241.585 43.985 ;
  END
 END o19
 PIN o20
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 43.795 240.825 44.365 ;
  END
 END o20
 PIN o21
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 44.175 241.585 44.745 ;
  END
 END o21
 PIN o22
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 44.555 240.825 45.125 ;
  END
 END o22
 PIN o23
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 44.935 241.585 45.505 ;
  END
 END o23
 PIN o24
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 45.315 240.825 45.885 ;
  END
 END o24
 PIN o25
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 45.695 241.585 46.265 ;
  END
 END o25
 PIN o26
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 46.075 240.825 46.645 ;
  END
 END o26
 PIN o27
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 47.215 241.585 47.785 ;
  END
 END o27
 PIN o28
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 47.595 240.825 48.165 ;
  END
 END o28
 PIN o29
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 47.975 241.585 48.545 ;
  END
 END o29
 PIN o30
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 49.495 241.585 50.065 ;
  END
 END o30
 PIN o31
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 49.875 240.825 50.445 ;
  END
 END o31
 PIN o32
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 50.255 241.585 50.825 ;
  END
 END o32
 PIN o33
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 68.115 241.585 68.685 ;
  END
 END o33
 PIN o34
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 68.875 241.585 69.445 ;
  END
 END o34
 PIN o35
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 70.395 241.585 70.965 ;
  END
 END o35
 PIN o36
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 70.775 240.825 71.345 ;
  END
 END o36
 PIN o37
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 71.155 241.585 71.725 ;
  END
 END o37
 PIN o38
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 71.535 240.825 72.105 ;
  END
 END o38
 PIN o39
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 50.635 240.825 51.205 ;
  END
 END o39
 PIN o40
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 52.535 241.585 53.105 ;
  END
 END o40
 PIN o41
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 52.915 240.825 53.485 ;
  END
 END o41
 PIN o42
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 53.675 241.585 54.245 ;
  END
 END o42
 PIN o43
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 54.055 240.825 54.625 ;
  END
 END o43
 PIN o44
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 54.435 241.585 55.005 ;
  END
 END o44
 PIN o45
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 54.815 240.825 55.385 ;
  END
 END o45
 PIN o46
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 55.195 241.585 55.765 ;
  END
 END o46
 PIN o47
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 56.335 241.585 56.905 ;
  END
 END o47
 PIN o48
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 56.715 240.825 57.285 ;
  END
 END o48
 PIN o49
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 57.095 241.585 57.665 ;
  END
 END o49
 PIN o50
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 57.475 240.825 58.045 ;
  END
 END o50
 PIN o51
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 57.855 241.585 58.425 ;
  END
 END o51
 PIN o52
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 58.235 240.825 58.805 ;
  END
 END o52
 PIN o53
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 58.615 241.585 59.185 ;
  END
 END o53
 PIN o54
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 58.995 240.825 59.565 ;
  END
 END o54
 PIN o55
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 59.375 241.585 59.945 ;
  END
 END o55
 PIN o56
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 59.755 240.825 60.325 ;
  END
 END o56
 PIN o57
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 63.935 124.545 64.505 125.115 ;
  END
 END o57
 PIN o58
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 67.355 124.545 67.925 125.115 ;
  END
 END o58
 PIN o59
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 80.655 124.545 81.225 125.115 ;
  END
 END o59
 PIN o60
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 98.515 124.545 99.085 125.115 ;
  END
 END o60
 PIN o61
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 48.355 3.325 48.925 ;
  END
 END o61
 PIN o62
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 40.375 3.325 40.945 ;
  END
 END o62
 PIN o63
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 39.615 3.325 40.185 ;
  END
 END o63
 PIN o64
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 47.975 4.085 48.545 ;
  END
 END o64
 PIN o65
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 44.935 3.325 45.505 ;
  END
 END o65
 PIN o66
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 44.175 3.325 44.745 ;
  END
 END o66
 PIN o67
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 124.545 130.245 125.115 ;
  END
 END o67
 PIN o68
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 135.375 124.545 135.945 125.115 ;
  END
 END o68
 PIN o69
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 168.435 124.545 169.005 125.115 ;
  END
 END o69
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 37.335 124.545 37.905 125.115 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 33.915 124.545 34.485 125.115 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 36.195 124.545 36.765 125.115 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 43.795 124.545 44.365 125.115 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 51.775 124.545 52.345 125.115 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 52.915 124.545 53.485 125.115 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 54.815 124.545 55.385 125.115 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 56.335 124.545 56.905 125.115 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 57.475 124.545 58.045 125.115 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 59.375 124.545 59.945 125.115 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 60.515 124.545 61.085 125.115 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 47.215 124.545 47.785 125.115 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 49.495 124.545 50.065 125.115 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 48.355 124.545 48.925 125.115 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 65.075 124.545 65.645 125.115 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 96.235 124.545 96.805 125.115 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 127.395 124.545 127.965 125.115 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 166.155 124.545 166.725 125.115 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 60.895 241.585 61.465 ;
  END
 END i18
 PIN i19
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 63.935 241.585 64.505 ;
  END
 END i19
 PIN i20
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 63.935 3.325 64.505 ;
  END
 END i20
 OBS
  LAYER metal1 ;
   RECT 0 0 244.72 126.54 ;
  LAYER via1 ;
   RECT 0 0 244.72 126.54 ;
  LAYER metal2 ;
   RECT 0 0 244.72 126.54 ;
  LAYER via2 ;
   RECT 0 0 244.72 126.54 ;
  LAYER metal3 ;
   RECT 0 0 244.72 126.54 ;
  LAYER via3 ;
   RECT 0 0 244.72 126.54 ;
  LAYER metal4 ;
   RECT 0 0 244.72 126.54 ;
 END
END block_644x666_91

MACRO block_321x324_66
 CLASS BLOCK ;
 FOREIGN block_321x324_66 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 121.98 BY 61.56 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 44.175 118.845 44.745 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 34.295 3.325 34.865 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 35.815 3.325 36.385 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 38.095 3.325 38.665 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 39.615 3.325 40.185 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 41.135 3.325 41.705 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 42.655 3.325 43.225 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 44.175 3.325 44.745 ;
  END
 END o7
 PIN o8
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 45.695 3.325 46.265 ;
  END
 END o8
 PIN o9
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 22.895 118.845 23.465 ;
  END
 END o9
 PIN o10
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 6.935 3.325 7.505 ;
  END
 END o10
 PIN o11
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 7.695 3.325 8.265 ;
  END
 END o11
 PIN o12
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 19.855 3.325 20.425 ;
  END
 END o12
 PIN o13
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 21.375 3.325 21.945 ;
  END
 END o13
 PIN o14
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 22.135 3.325 22.705 ;
  END
 END o14
 PIN o15
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 24.415 3.325 24.985 ;
  END
 END o15
 PIN o16
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 25.935 3.325 26.505 ;
  END
 END o16
 PIN o17
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 26.695 3.325 27.265 ;
  END
 END o17
 PIN o18
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 27.455 3.325 28.025 ;
  END
 END o18
 PIN o19
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 28.975 3.325 29.545 ;
  END
 END o19
 PIN o20
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 30.495 3.325 31.065 ;
  END
 END o20
 PIN o21
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 32.015 3.325 32.585 ;
  END
 END o21
 PIN o22
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 9.215 3.325 9.785 ;
  END
 END o22
 PIN o23
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 10.735 3.325 11.305 ;
  END
 END o23
 PIN o24
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 11.495 3.325 12.065 ;
  END
 END o24
 PIN o25
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 12.255 3.325 12.825 ;
  END
 END o25
 PIN o26
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 13.775 3.325 14.345 ;
  END
 END o26
 PIN o27
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 15.295 3.325 15.865 ;
  END
 END o27
 PIN o28
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 16.055 3.325 16.625 ;
  END
 END o28
 PIN o29
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 16.815 3.325 17.385 ;
  END
 END o29
 PIN o30
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 25.175 118.845 25.745 ;
  END
 END o30
 PIN o31
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 48.735 3.325 49.305 ;
  END
 END o31
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 32.015 118.845 32.585 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 44.935 118.845 45.505 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 30.495 118.845 31.065 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 31.255 118.845 31.825 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 35.055 118.845 35.625 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 34.295 118.845 34.865 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 27.455 118.845 28.025 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 28.975 118.845 29.545 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 24.415 118.845 24.985 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 42.655 118.845 43.225 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 47.215 3.325 47.785 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 4.655 3.325 5.225 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 22.135 118.845 22.705 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 21.375 118.845 21.945 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 29.735 118.845 30.305 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 26.695 118.845 27.265 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 25.935 118.845 26.505 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 3.895 118.845 4.465 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 4.655 118.845 5.225 ;
  END
 END i18
 PIN i19
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 6.175 118.845 6.745 ;
  END
 END i19
 PIN i20
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 6.935 118.845 7.505 ;
  END
 END i20
 PIN i21
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 7.695 118.845 8.265 ;
  END
 END i21
 PIN i22
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 8.455 118.845 9.025 ;
  END
 END i22
 PIN i23
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 9.215 118.845 9.785 ;
  END
 END i23
 PIN i24
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 10.735 118.845 11.305 ;
  END
 END i24
 PIN i25
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 11.495 118.845 12.065 ;
  END
 END i25
 PIN i26
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 12.255 118.845 12.825 ;
  END
 END i26
 PIN i27
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 13.015 118.845 13.585 ;
  END
 END i27
 PIN i28
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 13.775 118.845 14.345 ;
  END
 END i28
 PIN i29
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 15.295 118.845 15.865 ;
  END
 END i29
 PIN i30
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 16.055 118.845 16.625 ;
  END
 END i30
 PIN i31
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 16.815 118.845 17.385 ;
  END
 END i31
 PIN i32
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 17.575 118.845 18.145 ;
  END
 END i32
 PIN i33
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 18.335 118.845 18.905 ;
  END
 END i33
 OBS
  LAYER metal1 ;
   RECT 0 0 121.98 61.56 ;
  LAYER via1 ;
   RECT 0 0 121.98 61.56 ;
  LAYER metal2 ;
   RECT 0 0 121.98 61.56 ;
  LAYER via2 ;
   RECT 0 0 121.98 61.56 ;
  LAYER metal3 ;
   RECT 0 0 121.98 61.56 ;
  LAYER via3 ;
   RECT 0 0 121.98 61.56 ;
  LAYER metal4 ;
   RECT 0 0 121.98 61.56 ;
 END
END block_321x324_66

MACRO block_315x1863_130
 CLASS BLOCK ;
 FOREIGN block_315x1863_130 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 119.7 BY 353.97 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 298.395 9.785 298.965 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 304.095 9.785 304.665 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 315.685 9.785 316.255 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 321.385 9.785 321.955 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 2.565 9.785 3.135 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 19.665 9.785 20.235 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 25.555 9.785 26.125 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 31.255 9.785 31.825 ;
  END
 END o7
 PIN o8
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 36.955 9.785 37.525 ;
  END
 END o8
 PIN o9
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 327.085 9.785 327.655 ;
  END
 END o9
 PIN o10
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 48.545 9.785 49.115 ;
  END
 END o10
 PIN o11
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 54.245 9.785 54.815 ;
  END
 END o11
 PIN o12
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 59.945 9.785 60.515 ;
  END
 END o12
 PIN o13
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 71.535 9.785 72.105 ;
  END
 END o13
 PIN o14
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 77.235 9.785 77.805 ;
  END
 END o14
 PIN o15
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 82.935 9.785 83.505 ;
  END
 END o15
 PIN o16
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 88.635 9.785 89.205 ;
  END
 END o16
 PIN o17
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 94.525 9.785 95.095 ;
  END
 END o17
 PIN o18
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 100.225 9.785 100.795 ;
  END
 END o18
 PIN o19
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 105.925 9.785 106.495 ;
  END
 END o19
 PIN o20
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 128.915 9.785 129.485 ;
  END
 END o20
 PIN o21
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 134.615 9.785 135.185 ;
  END
 END o21
 PIN o22
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 140.505 9.785 141.075 ;
  END
 END o22
 PIN o23
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 151.905 9.785 152.475 ;
  END
 END o23
 PIN o24
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 338.675 9.785 339.245 ;
  END
 END o24
 PIN o25
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 157.605 9.785 158.175 ;
  END
 END o25
 PIN o26
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 163.495 9.785 164.065 ;
  END
 END o26
 PIN o27
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 212.135 9.785 212.705 ;
  END
 END o27
 PIN o28
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 223.725 9.785 224.295 ;
  END
 END o28
 PIN o29
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 235.125 9.785 235.695 ;
  END
 END o29
 PIN o30
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 241.015 9.785 241.585 ;
  END
 END o30
 PIN o31
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 246.715 9.785 247.285 ;
  END
 END o31
 PIN o32
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 252.415 9.785 252.985 ;
  END
 END o32
 PIN o33
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 258.115 9.785 258.685 ;
  END
 END o33
 PIN o34
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 264.005 9.785 264.575 ;
  END
 END o34
 PIN o35
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 269.705 9.785 270.275 ;
  END
 END o35
 PIN o36
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 281.105 9.785 281.675 ;
  END
 END o36
 PIN o37
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 286.995 9.785 287.565 ;
  END
 END o37
 PIN o38
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 292.695 9.785 293.265 ;
  END
 END o38
 PIN o39
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 344.375 9.785 344.945 ;
  END
 END o39
 PIN o40
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 350.075 9.785 350.645 ;
  END
 END o40
 PIN o41
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 65.645 9.785 66.215 ;
  END
 END o41
 PIN o42
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 275.405 9.785 275.975 ;
  END
 END o42
 PIN o43
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 195.035 9.785 195.605 ;
  END
 END o43
 PIN o44
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 200.735 9.785 201.305 ;
  END
 END o44
 PIN o45
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 123.215 9.785 123.785 ;
  END
 END o45
 PIN o46
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 218.025 9.785 218.595 ;
  END
 END o46
 PIN o47
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 206.435 9.785 207.005 ;
  END
 END o47
 PIN o48
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 332.975 9.785 333.545 ;
  END
 END o48
 PIN o49
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 309.985 9.785 310.555 ;
  END
 END o49
 PIN o50
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 229.425 9.785 229.995 ;
  END
 END o50
 PIN o51
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 146.205 9.785 146.775 ;
  END
 END o51
 PIN o52
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 111.625 9.785 112.195 ;
  END
 END o52
 PIN o53
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 117.515 9.785 118.085 ;
  END
 END o53
 PIN o54
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 42.655 9.785 43.225 ;
  END
 END o54
 PIN o55
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 8.265 9.785 8.835 ;
  END
 END o55
 PIN o56
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 13.965 9.785 14.535 ;
  END
 END o56
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 180.595 118.465 181.165 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 174.515 118.465 175.085 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 171.095 118.465 171.665 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.135 173.945 117.705 174.515 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 111.815 171.285 112.385 171.855 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 172.425 118.465 172.995 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 172.045 9.785 172.615 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 188.005 118.465 188.575 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 177.935 118.465 178.505 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 179.265 118.465 179.835 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 179.075 9.785 179.645 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 8.455 185.725 9.025 186.295 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 182.685 9.785 183.255 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.135 180.975 117.705 181.545 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 182.875 118.465 183.445 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.135 183.255 117.705 183.825 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 349.695 118.465 350.265 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 292.315 118.465 292.885 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 286.425 118.465 286.995 ;
  END
 END i18
 PIN i19
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 280.725 118.465 281.295 ;
  END
 END i19
 PIN i20
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 275.025 118.465 275.595 ;
  END
 END i20
 PIN i21
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 269.325 118.465 269.895 ;
  END
 END i21
 PIN i22
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 263.435 118.465 264.005 ;
  END
 END i22
 PIN i23
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 257.735 118.465 258.305 ;
  END
 END i23
 PIN i24
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 252.035 118.465 252.605 ;
  END
 END i24
 PIN i25
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 246.335 118.465 246.905 ;
  END
 END i25
 PIN i26
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 240.445 118.465 241.015 ;
  END
 END i26
 PIN i27
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 343.995 118.465 344.565 ;
  END
 END i27
 PIN i28
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 234.745 118.465 235.315 ;
  END
 END i28
 PIN i29
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 229.045 118.465 229.615 ;
  END
 END i29
 PIN i30
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 223.345 118.465 223.915 ;
  END
 END i30
 PIN i31
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 217.455 118.465 218.025 ;
  END
 END i31
 PIN i32
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 211.755 118.465 212.325 ;
  END
 END i32
 PIN i33
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 206.055 118.465 206.625 ;
  END
 END i33
 PIN i34
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 200.355 118.465 200.925 ;
  END
 END i34
 PIN i35
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 194.465 118.465 195.035 ;
  END
 END i35
 PIN i36
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 163.875 118.465 164.445 ;
  END
 END i36
 PIN i37
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 158.175 118.465 158.745 ;
  END
 END i37
 PIN i38
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 338.295 118.465 338.865 ;
  END
 END i38
 PIN i39
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 152.285 118.465 152.855 ;
  END
 END i39
 PIN i40
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 146.585 118.465 147.155 ;
  END
 END i40
 PIN i41
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 140.885 118.465 141.455 ;
  END
 END i41
 PIN i42
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 135.185 118.465 135.755 ;
  END
 END i42
 PIN i43
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 129.295 118.465 129.865 ;
  END
 END i43
 PIN i44
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 123.595 118.465 124.165 ;
  END
 END i44
 PIN i45
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 117.895 118.465 118.465 ;
  END
 END i45
 PIN i46
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 112.195 118.465 112.765 ;
  END
 END i46
 PIN i47
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 106.305 118.465 106.875 ;
  END
 END i47
 PIN i48
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 100.605 118.465 101.175 ;
  END
 END i48
 PIN i49
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 332.405 118.465 332.975 ;
  END
 END i49
 PIN i50
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 94.905 118.465 95.475 ;
  END
 END i50
 PIN i51
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 89.205 118.465 89.775 ;
  END
 END i51
 PIN i52
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 83.315 118.465 83.885 ;
  END
 END i52
 PIN i53
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 77.615 118.465 78.185 ;
  END
 END i53
 PIN i54
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 71.915 118.465 72.485 ;
  END
 END i54
 PIN i55
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 66.215 118.465 66.785 ;
  END
 END i55
 PIN i56
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 60.325 118.465 60.895 ;
  END
 END i56
 PIN i57
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 54.625 118.465 55.195 ;
  END
 END i57
 PIN i58
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 48.925 118.465 49.495 ;
  END
 END i58
 PIN i59
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 43.225 118.465 43.795 ;
  END
 END i59
 PIN i60
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 326.705 118.465 327.275 ;
  END
 END i60
 PIN i61
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 37.335 118.465 37.905 ;
  END
 END i61
 PIN i62
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 31.635 118.465 32.205 ;
  END
 END i62
 PIN i63
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 25.935 118.465 26.505 ;
  END
 END i63
 PIN i64
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 20.235 118.465 20.805 ;
  END
 END i64
 PIN i65
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 14.345 118.465 14.915 ;
  END
 END i65
 PIN i66
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 8.645 118.465 9.215 ;
  END
 END i66
 PIN i67
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 2.945 118.465 3.515 ;
  END
 END i67
 PIN i68
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 321.005 118.465 321.575 ;
  END
 END i68
 PIN i69
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 315.305 118.465 315.875 ;
  END
 END i69
 PIN i70
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 309.415 118.465 309.985 ;
  END
 END i70
 PIN i71
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 303.715 118.465 304.285 ;
  END
 END i71
 PIN i72
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 298.015 118.465 298.585 ;
  END
 END i72
 OBS
  LAYER metal1 ;
   RECT 0 0 119.7 353.97 ;
  LAYER via1 ;
   RECT 0 0 119.7 353.97 ;
  LAYER metal2 ;
   RECT 0 0 119.7 353.97 ;
  LAYER via2 ;
   RECT 0 0 119.7 353.97 ;
  LAYER metal3 ;
   RECT 0 0 119.7 353.97 ;
  LAYER via3 ;
   RECT 0 0 119.7 353.97 ;
  LAYER metal4 ;
   RECT 0 0 119.7 353.97 ;
 END
END block_315x1863_130

MACRO block_96x2070_138
 CLASS BLOCK ;
 FOREIGN block_96x2070_138 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 36.48 BY 393.3 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 19.855 9.785 20.425 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 25.555 9.785 26.125 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 59.945 9.785 60.515 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 65.835 9.785 66.405 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 100.225 9.785 100.795 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 105.925 9.785 106.495 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 88.825 9.785 89.395 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 128.915 9.785 129.485 ;
  END
 END o7
 PIN o8
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 111.815 9.785 112.385 ;
  END
 END o8
 PIN o9
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 31.255 9.785 31.825 ;
  END
 END o9
 PIN o10
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 71.535 9.785 72.105 ;
  END
 END o10
 PIN o11
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 212.325 9.785 212.895 ;
  END
 END o11
 PIN o12
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 146.205 9.785 146.775 ;
  END
 END o12
 PIN o13
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 252.415 9.785 252.985 ;
  END
 END o13
 PIN o14
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 292.695 9.785 293.265 ;
  END
 END o14
 PIN o15
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 140.505 9.785 141.075 ;
  END
 END o15
 PIN o16
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 246.715 9.785 247.285 ;
  END
 END o16
 PIN o17
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 180.785 9.785 181.355 ;
  END
 END o17
 PIN o18
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 286.995 9.785 287.565 ;
  END
 END o18
 PIN o19
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 117.515 9.785 118.085 ;
  END
 END o19
 PIN o20
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 298.395 9.785 298.965 ;
  END
 END o20
 PIN o21
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 77.235 9.785 77.805 ;
  END
 END o21
 PIN o22
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 36.955 9.785 37.525 ;
  END
 END o22
 PIN o23
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 258.305 9.785 258.875 ;
  END
 END o23
 PIN o24
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 218.025 9.785 218.595 ;
  END
 END o24
 PIN o25
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 327.275 9.785 327.845 ;
  END
 END o25
 PIN o26
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 361.665 9.785 362.235 ;
  END
 END o26
 PIN o27
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 378.955 9.785 379.525 ;
  END
 END o27
 PIN o28
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 344.375 9.785 344.945 ;
  END
 END o28
 PIN o29
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 223.725 9.785 224.295 ;
  END
 END o29
 PIN o30
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 264.005 9.785 264.575 ;
  END
 END o30
 PIN o31
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 304.285 9.785 304.855 ;
  END
 END o31
 PIN o32
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 275.405 9.785 275.975 ;
  END
 END o32
 PIN o33
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 315.685 9.785 316.255 ;
  END
 END o33
 PIN o34
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 350.265 9.785 350.835 ;
  END
 END o34
 PIN o35
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 269.705 9.785 270.275 ;
  END
 END o35
 PIN o36
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 229.425 9.785 229.995 ;
  END
 END o36
 PIN o37
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 384.655 9.785 385.225 ;
  END
 END o37
 PIN o38
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 235.315 9.785 235.885 ;
  END
 END o38
 PIN o39
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 48.545 9.785 49.115 ;
  END
 END o39
 PIN o40
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 8.265 9.785 8.835 ;
  END
 END o40
 PIN o41
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 54.245 9.785 54.815 ;
  END
 END o41
 PIN o42
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 367.365 9.785 367.935 ;
  END
 END o42
 PIN o43
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 373.255 9.785 373.825 ;
  END
 END o43
 PIN o44
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 390.355 9.785 390.925 ;
  END
 END o44
 PIN o45
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 332.975 9.785 333.545 ;
  END
 END o45
 PIN o46
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 338.675 9.785 339.245 ;
  END
 END o46
 PIN o47
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 309.985 9.785 310.555 ;
  END
 END o47
 PIN o48
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 151.905 9.785 152.475 ;
  END
 END o48
 PIN o49
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 157.795 9.785 158.365 ;
  END
 END o49
 PIN o50
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 169.195 9.785 169.765 ;
  END
 END o50
 PIN o51
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 163.495 9.785 164.065 ;
  END
 END o51
 PIN o52
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 123.215 9.785 123.785 ;
  END
 END o52
 PIN o53
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 134.805 9.785 135.375 ;
  END
 END o53
 PIN o54
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 82.935 9.785 83.505 ;
  END
 END o54
 PIN o55
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 94.525 9.785 95.095 ;
  END
 END o55
 PIN o56
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 42.845 9.785 43.415 ;
  END
 END o56
 PIN o57
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 2.565 9.785 3.135 ;
  END
 END o57
 PIN o58
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 13.965 9.785 14.535 ;
  END
 END o58
 PIN o59
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 174.895 9.785 175.465 ;
  END
 END o59
 PIN o60
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 355.965 9.785 356.535 ;
  END
 END o60
 PIN o61
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 321.385 9.785 321.955 ;
  END
 END o61
 PIN o62
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 281.295 9.785 281.865 ;
  END
 END o62
 PIN o63
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 241.015 9.785 241.585 ;
  END
 END o63
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 197.885 35.245 198.455 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 188.385 35.245 188.955 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 188.575 29.165 189.145 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 189.335 9.785 189.905 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 205.295 35.245 205.865 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 195.225 35.245 195.795 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 196.555 35.245 197.125 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 196.365 9.785 196.935 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 8.455 203.015 9.025 203.585 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 199.975 9.785 200.545 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 389.975 35.245 390.545 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 332.595 35.245 333.165 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 326.705 35.245 327.275 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 321.005 35.245 321.575 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 315.305 35.245 315.875 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 309.605 35.245 310.175 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 303.715 35.245 304.285 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 298.015 35.245 298.585 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 292.315 35.245 292.885 ;
  END
 END i18
 PIN i19
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 286.615 35.245 287.185 ;
  END
 END i19
 PIN i20
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 280.725 35.245 281.295 ;
  END
 END i20
 PIN i21
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 384.275 35.245 384.845 ;
  END
 END i21
 PIN i22
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 275.025 35.245 275.595 ;
  END
 END i22
 PIN i23
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 269.325 35.245 269.895 ;
  END
 END i23
 PIN i24
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 263.625 35.245 264.195 ;
  END
 END i24
 PIN i25
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 257.735 35.245 258.305 ;
  END
 END i25
 PIN i26
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 252.035 35.245 252.605 ;
  END
 END i26
 PIN i27
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 246.335 35.245 246.905 ;
  END
 END i27
 PIN i28
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 240.635 35.245 241.205 ;
  END
 END i28
 PIN i29
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 234.745 35.245 235.315 ;
  END
 END i29
 PIN i30
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 229.045 35.245 229.615 ;
  END
 END i30
 PIN i31
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 223.345 35.245 223.915 ;
  END
 END i31
 PIN i32
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 378.575 35.245 379.145 ;
  END
 END i32
 PIN i33
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 217.645 35.245 218.215 ;
  END
 END i33
 PIN i34
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 211.755 35.245 212.325 ;
  END
 END i34
 PIN i35
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 181.165 35.245 181.735 ;
  END
 END i35
 PIN i36
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 175.465 35.245 176.035 ;
  END
 END i36
 PIN i37
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 169.575 35.245 170.145 ;
  END
 END i37
 PIN i38
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 163.875 35.245 164.445 ;
  END
 END i38
 PIN i39
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 158.175 35.245 158.745 ;
  END
 END i39
 PIN i40
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 152.475 35.245 153.045 ;
  END
 END i40
 PIN i41
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 146.585 35.245 147.155 ;
  END
 END i41
 PIN i42
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 140.885 35.245 141.455 ;
  END
 END i42
 PIN i43
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 372.685 35.245 373.255 ;
  END
 END i43
 PIN i44
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 135.185 35.245 135.755 ;
  END
 END i44
 PIN i45
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 129.485 35.245 130.055 ;
  END
 END i45
 PIN i46
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 123.595 35.245 124.165 ;
  END
 END i46
 PIN i47
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 117.895 35.245 118.465 ;
  END
 END i47
 PIN i48
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 112.195 35.245 112.765 ;
  END
 END i48
 PIN i49
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 106.495 35.245 107.065 ;
  END
 END i49
 PIN i50
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 100.605 35.245 101.175 ;
  END
 END i50
 PIN i51
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 94.905 35.245 95.475 ;
  END
 END i51
 PIN i52
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 89.205 35.245 89.775 ;
  END
 END i52
 PIN i53
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 83.505 35.245 84.075 ;
  END
 END i53
 PIN i54
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 366.985 35.245 367.555 ;
  END
 END i54
 PIN i55
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 77.615 35.245 78.185 ;
  END
 END i55
 PIN i56
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 71.915 35.245 72.485 ;
  END
 END i56
 PIN i57
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 66.215 35.245 66.785 ;
  END
 END i57
 PIN i58
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 60.515 35.245 61.085 ;
  END
 END i58
 PIN i59
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 54.625 35.245 55.195 ;
  END
 END i59
 PIN i60
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 48.925 35.245 49.495 ;
  END
 END i60
 PIN i61
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 43.225 35.245 43.795 ;
  END
 END i61
 PIN i62
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 37.525 35.245 38.095 ;
  END
 END i62
 PIN i63
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 31.635 35.245 32.205 ;
  END
 END i63
 PIN i64
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 25.935 35.245 26.505 ;
  END
 END i64
 PIN i65
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 361.285 35.245 361.855 ;
  END
 END i65
 PIN i66
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 20.235 35.245 20.805 ;
  END
 END i66
 PIN i67
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 14.535 35.245 15.105 ;
  END
 END i67
 PIN i68
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 8.645 35.245 9.215 ;
  END
 END i68
 PIN i69
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 2.945 35.245 3.515 ;
  END
 END i69
 PIN i70
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 355.585 35.245 356.155 ;
  END
 END i70
 PIN i71
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 349.695 35.245 350.265 ;
  END
 END i71
 PIN i72
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 343.995 35.245 344.565 ;
  END
 END i72
 PIN i73
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.675 338.295 35.245 338.865 ;
  END
 END i73
 OBS
  LAYER metal1 ;
   RECT 0 0 36.48 393.3 ;
  LAYER via1 ;
   RECT 0 0 36.48 393.3 ;
  LAYER metal2 ;
   RECT 0 0 36.48 393.3 ;
  LAYER via2 ;
   RECT 0 0 36.48 393.3 ;
  LAYER metal3 ;
   RECT 0 0 36.48 393.3 ;
  LAYER via3 ;
   RECT 0 0 36.48 393.3 ;
  LAYER metal4 ;
   RECT 0 0 36.48 393.3 ;
 END
END block_96x2070_138

MACRO block_737x3078_1192
 CLASS BLOCK ;
 FOREIGN block_737x3078_1192 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 280.06 BY 584.82 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 582.255 268.565 582.825 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 255.835 582.255 256.405 582.825 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 237.975 582.255 238.545 582.825 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 239.115 582.255 239.685 582.825 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 236.075 582.255 236.645 582.825 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 139.555 582.255 140.125 582.825 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 138.415 582.255 138.985 582.825 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 136.515 582.255 137.085 582.825 ;
  END
 END o7
 PIN o8
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 145.635 582.255 146.205 582.825 ;
  END
 END o8
 PIN o9
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 144.495 582.255 145.065 582.825 ;
  END
 END o9
 PIN o10
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 170.335 582.255 170.905 582.825 ;
  END
 END o10
 PIN o11
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 226.955 582.255 227.525 582.825 ;
  END
 END o11
 PIN o12
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 225.815 582.255 226.385 582.825 ;
  END
 END o12
 PIN o13
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 223.915 582.255 224.485 582.825 ;
  END
 END o13
 PIN o14
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 233.035 582.255 233.605 582.825 ;
  END
 END o14
 PIN o15
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 153.615 582.255 154.185 582.825 ;
  END
 END o15
 PIN o16
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 151.715 582.255 152.285 582.825 ;
  END
 END o16
 PIN o17
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 150.575 582.255 151.145 582.825 ;
  END
 END o17
 PIN o18
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 252.795 582.255 253.365 582.825 ;
  END
 END o18
 PIN o19
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 251.655 582.255 252.225 582.825 ;
  END
 END o19
 PIN o20
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.515 582.255 175.085 582.825 ;
  END
 END o20
 PIN o21
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 171.475 582.255 172.045 582.825 ;
  END
 END o21
 PIN o22
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 173.375 582.255 173.945 582.825 ;
  END
 END o22
 PIN o23
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 231.895 582.255 232.465 582.825 ;
  END
 END o23
 PIN o24
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 234.935 582.255 235.505 582.825 ;
  END
 END o24
 PIN o25
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 147.535 582.255 148.105 582.825 ;
  END
 END o25
 PIN o26
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 148.675 582.255 149.245 582.825 ;
  END
 END o26
 PIN o27
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.755 582.255 155.325 582.825 ;
  END
 END o27
 PIN o28
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 157.795 582.255 158.365 582.825 ;
  END
 END o28
 PIN o29
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 159.695 582.255 160.265 582.825 ;
  END
 END o29
 PIN o30
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 182.495 582.255 183.065 582.825 ;
  END
 END o30
 PIN o31
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 183.635 582.255 184.205 582.825 ;
  END
 END o31
 PIN o32
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 185.535 582.255 186.105 582.825 ;
  END
 END o32
 PIN o33
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 180.595 582.255 181.165 582.825 ;
  END
 END o33
 PIN o34
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 177.555 582.255 178.125 582.825 ;
  END
 END o34
 PIN o35
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.895 582.255 270.465 582.825 ;
  END
 END o35
 PIN o36
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 258.875 582.255 259.445 582.825 ;
  END
 END o36
 PIN o37
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 271.035 582.255 271.605 582.825 ;
  END
 END o37
 PIN o38
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 245.195 582.255 245.765 582.825 ;
  END
 END o38
 PIN o39
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 165.395 582.255 165.965 582.825 ;
  END
 END o39
 PIN o40
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 162.355 582.255 162.925 582.825 ;
  END
 END o40
 PIN o41
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 249.755 582.255 250.325 582.825 ;
  END
 END o41
 PIN o42
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 261.915 582.255 262.485 582.825 ;
  END
 END o42
 PIN o43
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 247.095 582.255 247.665 582.825 ;
  END
 END o43
 PIN o44
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 263.815 582.255 264.385 582.825 ;
  END
 END o44
 PIN o45
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 264.955 582.255 265.525 582.825 ;
  END
 END o45
 PIN o46
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 266.855 582.255 267.425 582.825 ;
  END
 END o46
 PIN o47
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 168.435 582.255 169.005 582.825 ;
  END
 END o47
 PIN o48
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 176.415 582.255 176.985 582.825 ;
  END
 END o48
 PIN o49
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 179.455 582.255 180.025 582.825 ;
  END
 END o49
 PIN o50
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 257.735 582.255 258.305 582.825 ;
  END
 END o50
 PIN o51
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 260.775 582.255 261.345 582.825 ;
  END
 END o51
 PIN o52
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 254.695 582.255 255.265 582.825 ;
  END
 END o52
 PIN o53
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 142.595 582.255 143.165 582.825 ;
  END
 END o53
 PIN o54
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 229.995 582.255 230.565 582.825 ;
  END
 END o54
 PIN o55
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 228.855 582.255 229.425 582.825 ;
  END
 END o55
 PIN o56
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 582.255 241.585 582.825 ;
  END
 END o56
 PIN o57
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 167.295 582.255 167.865 582.825 ;
  END
 END o57
 PIN o58
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 164.255 582.255 164.825 582.825 ;
  END
 END o58
 PIN o59
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 242.155 582.255 242.725 582.825 ;
  END
 END o59
 PIN o60
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 141.455 582.255 142.025 582.825 ;
  END
 END o60
 PIN o61
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 272.935 582.255 273.505 582.825 ;
  END
 END o61
 PIN o62
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 244.055 582.255 244.625 582.825 ;
  END
 END o62
 PIN o63
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 156.655 582.255 157.225 582.825 ;
  END
 END o63
 PIN o64
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 205.295 582.255 205.865 582.825 ;
  END
 END o64
 PIN o65
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.915 0.665 72.485 1.235 ;
  END
 END o65
 PIN o66
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 29.355 582.255 29.925 582.825 ;
  END
 END o66
 PIN o67
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 47.405 3.325 47.975 ;
  END
 END o67
 PIN o68
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 48.165 3.325 48.735 ;
  END
 END o68
 PIN o69
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 103.645 3.325 104.215 ;
  END
 END o69
 PIN o70
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 347.415 3.325 347.985 ;
  END
 END o70
 PIN o71
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 351.025 3.325 351.595 ;
  END
 END o71
 PIN o72
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 351.785 3.325 352.355 ;
  END
 END o72
 PIN o73
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 355.395 3.325 355.965 ;
  END
 END o73
 PIN o74
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 356.155 3.325 356.725 ;
  END
 END o74
 PIN o75
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 359.765 3.325 360.335 ;
  END
 END o75
 PIN o76
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 360.525 3.325 361.095 ;
  END
 END o76
 PIN o77
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 364.135 3.325 364.705 ;
  END
 END o77
 PIN o78
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 364.895 3.325 365.465 ;
  END
 END o78
 PIN o79
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 368.505 3.325 369.075 ;
  END
 END o79
 PIN o80
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 104.405 3.325 104.975 ;
  END
 END o80
 PIN o81
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 369.265 3.325 369.835 ;
  END
 END o81
 PIN o82
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 372.875 3.325 373.445 ;
  END
 END o82
 PIN o83
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 373.635 3.325 374.205 ;
  END
 END o83
 PIN o84
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 377.245 3.325 377.815 ;
  END
 END o84
 PIN o85
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 378.005 3.325 378.575 ;
  END
 END o85
 PIN o86
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 381.615 3.325 382.185 ;
  END
 END o86
 PIN o87
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 382.375 3.325 382.945 ;
  END
 END o87
 PIN o88
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 385.985 3.325 386.555 ;
  END
 END o88
 PIN o89
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 402.135 3.325 402.705 ;
  END
 END o89
 PIN o90
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 402.895 3.325 403.465 ;
  END
 END o90
 PIN o91
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 108.015 3.325 108.585 ;
  END
 END o91
 PIN o92
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 440.895 3.325 441.465 ;
  END
 END o92
 PIN o93
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 441.655 3.325 442.225 ;
  END
 END o93
 PIN o94
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 445.265 3.325 445.835 ;
  END
 END o94
 PIN o95
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 446.025 3.325 446.595 ;
  END
 END o95
 PIN o96
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 449.635 3.325 450.205 ;
  END
 END o96
 PIN o97
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 450.395 3.325 450.965 ;
  END
 END o97
 PIN o98
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 454.005 3.325 454.575 ;
  END
 END o98
 PIN o99
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 454.765 3.325 455.335 ;
  END
 END o99
 PIN o100
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 458.375 3.325 458.945 ;
  END
 END o100
 PIN o101
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 459.135 3.325 459.705 ;
  END
 END o101
 PIN o102
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 108.775 3.325 109.345 ;
  END
 END o102
 PIN o103
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 462.745 3.325 463.315 ;
  END
 END o103
 PIN o104
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 463.505 3.325 464.075 ;
  END
 END o104
 PIN o105
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 467.115 3.325 467.685 ;
  END
 END o105
 PIN o106
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 467.875 3.325 468.445 ;
  END
 END o106
 PIN o107
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 471.485 3.325 472.055 ;
  END
 END o107
 PIN o108
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 472.245 3.325 472.815 ;
  END
 END o108
 PIN o109
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 475.855 3.325 476.425 ;
  END
 END o109
 PIN o110
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 476.615 3.325 477.185 ;
  END
 END o110
 PIN o111
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 480.225 3.325 480.795 ;
  END
 END o111
 PIN o112
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 480.985 3.325 481.555 ;
  END
 END o112
 PIN o113
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 112.385 3.325 112.955 ;
  END
 END o113
 PIN o114
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 484.595 3.325 485.165 ;
  END
 END o114
 PIN o115
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 485.355 3.325 485.925 ;
  END
 END o115
 PIN o116
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 488.965 3.325 489.535 ;
  END
 END o116
 PIN o117
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 489.725 3.325 490.295 ;
  END
 END o117
 PIN o118
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 493.335 3.325 493.905 ;
  END
 END o118
 PIN o119
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 494.095 3.325 494.665 ;
  END
 END o119
 PIN o120
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 497.705 3.325 498.275 ;
  END
 END o120
 PIN o121
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 498.465 3.325 499.035 ;
  END
 END o121
 PIN o122
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 502.075 3.325 502.645 ;
  END
 END o122
 PIN o123
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 502.835 3.325 503.405 ;
  END
 END o123
 PIN o124
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 113.145 3.325 113.715 ;
  END
 END o124
 PIN o125
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 506.445 3.325 507.015 ;
  END
 END o125
 PIN o126
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 507.205 3.325 507.775 ;
  END
 END o126
 PIN o127
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 510.815 3.325 511.385 ;
  END
 END o127
 PIN o128
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 511.575 3.325 512.145 ;
  END
 END o128
 PIN o129
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 515.185 3.325 515.755 ;
  END
 END o129
 PIN o130
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 515.945 3.325 516.515 ;
  END
 END o130
 PIN o131
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 519.555 3.325 520.125 ;
  END
 END o131
 PIN o132
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 520.315 3.325 520.885 ;
  END
 END o132
 PIN o133
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 523.925 3.325 524.495 ;
  END
 END o133
 PIN o134
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 524.685 3.325 525.255 ;
  END
 END o134
 PIN o135
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 116.755 3.325 117.325 ;
  END
 END o135
 PIN o136
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 528.295 3.325 528.865 ;
  END
 END o136
 PIN o137
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 529.055 3.325 529.625 ;
  END
 END o137
 PIN o138
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 532.665 3.325 533.235 ;
  END
 END o138
 PIN o139
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 533.425 3.325 533.995 ;
  END
 END o139
 PIN o140
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 537.035 3.325 537.605 ;
  END
 END o140
 PIN o141
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 537.795 3.325 538.365 ;
  END
 END o141
 PIN o142
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 541.405 3.325 541.975 ;
  END
 END o142
 PIN o143
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 542.165 3.325 542.735 ;
  END
 END o143
 PIN o144
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 545.775 3.325 546.345 ;
  END
 END o144
 PIN o145
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 546.535 3.325 547.105 ;
  END
 END o145
 PIN o146
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 117.515 3.325 118.085 ;
  END
 END o146
 PIN o147
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 550.145 3.325 550.715 ;
  END
 END o147
 PIN o148
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 550.905 3.325 551.475 ;
  END
 END o148
 PIN o149
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 554.515 3.325 555.085 ;
  END
 END o149
 PIN o150
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 555.275 3.325 555.845 ;
  END
 END o150
 PIN o151
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 558.885 3.325 559.455 ;
  END
 END o151
 PIN o152
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 559.645 3.325 560.215 ;
  END
 END o152
 PIN o153
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 563.255 3.325 563.825 ;
  END
 END o153
 PIN o154
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 121.125 3.325 121.695 ;
  END
 END o154
 PIN o155
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 121.885 3.325 122.455 ;
  END
 END o155
 PIN o156
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 86.165 3.325 86.735 ;
  END
 END o156
 PIN o157
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 125.495 3.325 126.065 ;
  END
 END o157
 PIN o158
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 126.255 3.325 126.825 ;
  END
 END o158
 PIN o159
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 129.865 3.325 130.435 ;
  END
 END o159
 PIN o160
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 130.625 3.325 131.195 ;
  END
 END o160
 PIN o161
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 134.235 3.325 134.805 ;
  END
 END o161
 PIN o162
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 134.995 3.325 135.565 ;
  END
 END o162
 PIN o163
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 138.605 3.325 139.175 ;
  END
 END o163
 PIN o164
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 139.365 3.325 139.935 ;
  END
 END o164
 PIN o165
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 142.975 3.325 143.545 ;
  END
 END o165
 PIN o166
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 143.735 3.325 144.305 ;
  END
 END o166
 PIN o167
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 86.925 3.325 87.495 ;
  END
 END o167
 PIN o168
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 147.345 3.325 147.915 ;
  END
 END o168
 PIN o169
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 148.105 3.325 148.675 ;
  END
 END o169
 PIN o170
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 151.715 3.325 152.285 ;
  END
 END o170
 PIN o171
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 152.475 3.325 153.045 ;
  END
 END o171
 PIN o172
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 156.085 3.325 156.655 ;
  END
 END o172
 PIN o173
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 156.845 3.325 157.415 ;
  END
 END o173
 PIN o174
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 160.455 3.325 161.025 ;
  END
 END o174
 PIN o175
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 161.215 3.325 161.785 ;
  END
 END o175
 PIN o176
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 164.825 3.325 165.395 ;
  END
 END o176
 PIN o177
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 165.585 3.325 166.155 ;
  END
 END o177
 PIN o178
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 90.535 3.325 91.105 ;
  END
 END o178
 PIN o179
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 169.195 3.325 169.765 ;
  END
 END o179
 PIN o180
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 169.955 3.325 170.525 ;
  END
 END o180
 PIN o181
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 173.565 3.325 174.135 ;
  END
 END o181
 PIN o182
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 174.325 3.325 174.895 ;
  END
 END o182
 PIN o183
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 177.935 3.325 178.505 ;
  END
 END o183
 PIN o184
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 178.695 3.325 179.265 ;
  END
 END o184
 PIN o185
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 182.305 3.325 182.875 ;
  END
 END o185
 PIN o186
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 183.065 3.325 183.635 ;
  END
 END o186
 PIN o187
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 186.675 3.325 187.245 ;
  END
 END o187
 PIN o188
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 187.435 3.325 188.005 ;
  END
 END o188
 PIN o189
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 91.295 3.325 91.865 ;
  END
 END o189
 PIN o190
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 191.045 3.325 191.615 ;
  END
 END o190
 PIN o191
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 191.805 3.325 192.375 ;
  END
 END o191
 PIN o192
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 195.415 3.325 195.985 ;
  END
 END o192
 PIN o193
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 196.175 3.325 196.745 ;
  END
 END o193
 PIN o194
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 199.785 3.325 200.355 ;
  END
 END o194
 PIN o195
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 200.545 3.325 201.115 ;
  END
 END o195
 PIN o196
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 204.155 3.325 204.725 ;
  END
 END o196
 PIN o197
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 204.915 3.325 205.485 ;
  END
 END o197
 PIN o198
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 208.525 3.325 209.095 ;
  END
 END o198
 PIN o199
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 224.675 3.325 225.245 ;
  END
 END o199
 PIN o200
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 94.905 3.325 95.475 ;
  END
 END o200
 PIN o201
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 225.435 3.325 226.005 ;
  END
 END o201
 PIN o202
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 263.625 3.325 264.195 ;
  END
 END o202
 PIN o203
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 264.385 3.325 264.955 ;
  END
 END o203
 PIN o204
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 267.995 3.325 268.565 ;
  END
 END o204
 PIN o205
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 268.755 3.325 269.325 ;
  END
 END o205
 PIN o206
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 272.365 3.325 272.935 ;
  END
 END o206
 PIN o207
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 273.125 3.325 273.695 ;
  END
 END o207
 PIN o208
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 276.735 3.325 277.305 ;
  END
 END o208
 PIN o209
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 277.495 3.325 278.065 ;
  END
 END o209
 PIN o210
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 281.105 3.325 281.675 ;
  END
 END o210
 PIN o211
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 95.665 3.325 96.235 ;
  END
 END o211
 PIN o212
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 281.865 3.325 282.435 ;
  END
 END o212
 PIN o213
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 285.475 3.325 286.045 ;
  END
 END o213
 PIN o214
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 286.235 3.325 286.805 ;
  END
 END o214
 PIN o215
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 289.845 3.325 290.415 ;
  END
 END o215
 PIN o216
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 290.605 3.325 291.175 ;
  END
 END o216
 PIN o217
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 294.215 3.325 294.785 ;
  END
 END o217
 PIN o218
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 294.975 3.325 295.545 ;
  END
 END o218
 PIN o219
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 298.585 3.325 299.155 ;
  END
 END o219
 PIN o220
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 299.345 3.325 299.915 ;
  END
 END o220
 PIN o221
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 302.955 3.325 303.525 ;
  END
 END o221
 PIN o222
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 99.275 3.325 99.845 ;
  END
 END o222
 PIN o223
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 303.715 3.325 304.285 ;
  END
 END o223
 PIN o224
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 307.325 3.325 307.895 ;
  END
 END o224
 PIN o225
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 308.085 3.325 308.655 ;
  END
 END o225
 PIN o226
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 311.695 3.325 312.265 ;
  END
 END o226
 PIN o227
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 312.455 3.325 313.025 ;
  END
 END o227
 PIN o228
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 316.065 3.325 316.635 ;
  END
 END o228
 PIN o229
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 316.825 3.325 317.395 ;
  END
 END o229
 PIN o230
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 320.435 3.325 321.005 ;
  END
 END o230
 PIN o231
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 321.195 3.325 321.765 ;
  END
 END o231
 PIN o232
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 324.805 3.325 325.375 ;
  END
 END o232
 PIN o233
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 100.035 3.325 100.605 ;
  END
 END o233
 PIN o234
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 325.565 3.325 326.135 ;
  END
 END o234
 PIN o235
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 329.175 3.325 329.745 ;
  END
 END o235
 PIN o236
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 329.935 3.325 330.505 ;
  END
 END o236
 PIN o237
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 333.545 3.325 334.115 ;
  END
 END o237
 PIN o238
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 334.305 3.325 334.875 ;
  END
 END o238
 PIN o239
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 337.915 3.325 338.485 ;
  END
 END o239
 PIN o240
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 338.675 3.325 339.245 ;
  END
 END o240
 PIN o241
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 342.285 3.325 342.855 ;
  END
 END o241
 PIN o242
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 343.045 3.325 343.615 ;
  END
 END o242
 PIN o243
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 346.655 3.325 347.225 ;
  END
 END o243
 PIN o244
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 46.835 29.165 47.405 ;
  END
 END o244
 PIN o245
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 49.115 29.165 49.685 ;
  END
 END o245
 PIN o246
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 103.455 29.165 104.025 ;
  END
 END o246
 PIN o247
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 347.795 29.165 348.365 ;
  END
 END o247
 PIN o248
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 350.835 29.165 351.405 ;
  END
 END o248
 PIN o249
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 352.165 29.165 352.735 ;
  END
 END o249
 PIN o250
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 355.205 29.165 355.775 ;
  END
 END o250
 PIN o251
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 356.535 29.165 357.105 ;
  END
 END o251
 PIN o252
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 359.575 29.165 360.145 ;
  END
 END o252
 PIN o253
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 360.905 29.165 361.475 ;
  END
 END o253
 PIN o254
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 363.945 29.165 364.515 ;
  END
 END o254
 PIN o255
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 365.275 29.165 365.845 ;
  END
 END o255
 PIN o256
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 368.315 29.165 368.885 ;
  END
 END o256
 PIN o257
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 104.785 29.165 105.355 ;
  END
 END o257
 PIN o258
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 369.645 29.165 370.215 ;
  END
 END o258
 PIN o259
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 372.685 29.165 373.255 ;
  END
 END o259
 PIN o260
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 374.015 29.165 374.585 ;
  END
 END o260
 PIN o261
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 377.055 29.165 377.625 ;
  END
 END o261
 PIN o262
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 378.385 29.165 378.955 ;
  END
 END o262
 PIN o263
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 381.425 29.165 381.995 ;
  END
 END o263
 PIN o264
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 382.755 29.165 383.325 ;
  END
 END o264
 PIN o265
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 385.795 29.165 386.365 ;
  END
 END o265
 PIN o266
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 401.565 29.165 402.135 ;
  END
 END o266
 PIN o267
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 403.845 29.165 404.415 ;
  END
 END o267
 PIN o268
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 107.825 29.165 108.395 ;
  END
 END o268
 PIN o269
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 440.705 29.165 441.275 ;
  END
 END o269
 PIN o270
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 442.035 29.165 442.605 ;
  END
 END o270
 PIN o271
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 445.075 29.165 445.645 ;
  END
 END o271
 PIN o272
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 446.405 29.165 446.975 ;
  END
 END o272
 PIN o273
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 449.445 29.165 450.015 ;
  END
 END o273
 PIN o274
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 450.775 29.165 451.345 ;
  END
 END o274
 PIN o275
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 453.815 29.165 454.385 ;
  END
 END o275
 PIN o276
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 455.145 29.165 455.715 ;
  END
 END o276
 PIN o277
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 458.185 29.165 458.755 ;
  END
 END o277
 PIN o278
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 459.515 29.165 460.085 ;
  END
 END o278
 PIN o279
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 109.155 29.165 109.725 ;
  END
 END o279
 PIN o280
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 462.555 29.165 463.125 ;
  END
 END o280
 PIN o281
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 463.885 29.165 464.455 ;
  END
 END o281
 PIN o282
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 466.925 29.165 467.495 ;
  END
 END o282
 PIN o283
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 468.255 29.165 468.825 ;
  END
 END o283
 PIN o284
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 471.295 29.165 471.865 ;
  END
 END o284
 PIN o285
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 472.625 29.165 473.195 ;
  END
 END o285
 PIN o286
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 475.665 29.165 476.235 ;
  END
 END o286
 PIN o287
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 476.995 29.165 477.565 ;
  END
 END o287
 PIN o288
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 480.035 29.165 480.605 ;
  END
 END o288
 PIN o289
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 481.365 29.165 481.935 ;
  END
 END o289
 PIN o290
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 112.195 29.165 112.765 ;
  END
 END o290
 PIN o291
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 484.405 29.165 484.975 ;
  END
 END o291
 PIN o292
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 485.735 29.165 486.305 ;
  END
 END o292
 PIN o293
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 488.775 29.165 489.345 ;
  END
 END o293
 PIN o294
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 490.105 29.165 490.675 ;
  END
 END o294
 PIN o295
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 493.145 29.165 493.715 ;
  END
 END o295
 PIN o296
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 494.475 29.165 495.045 ;
  END
 END o296
 PIN o297
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 497.515 29.165 498.085 ;
  END
 END o297
 PIN o298
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 498.845 29.165 499.415 ;
  END
 END o298
 PIN o299
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 501.885 29.165 502.455 ;
  END
 END o299
 PIN o300
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 503.215 29.165 503.785 ;
  END
 END o300
 PIN o301
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 113.525 29.165 114.095 ;
  END
 END o301
 PIN o302
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 506.255 29.165 506.825 ;
  END
 END o302
 PIN o303
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 507.585 29.165 508.155 ;
  END
 END o303
 PIN o304
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 510.625 29.165 511.195 ;
  END
 END o304
 PIN o305
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 511.955 29.165 512.525 ;
  END
 END o305
 PIN o306
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 514.995 29.165 515.565 ;
  END
 END o306
 PIN o307
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 516.325 29.165 516.895 ;
  END
 END o307
 PIN o308
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 519.365 29.165 519.935 ;
  END
 END o308
 PIN o309
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 520.695 29.165 521.265 ;
  END
 END o309
 PIN o310
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 523.735 29.165 524.305 ;
  END
 END o310
 PIN o311
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 525.065 29.165 525.635 ;
  END
 END o311
 PIN o312
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 116.565 29.165 117.135 ;
  END
 END o312
 PIN o313
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 528.105 29.165 528.675 ;
  END
 END o313
 PIN o314
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 529.435 29.165 530.005 ;
  END
 END o314
 PIN o315
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 532.475 29.165 533.045 ;
  END
 END o315
 PIN o316
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 533.805 29.165 534.375 ;
  END
 END o316
 PIN o317
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 536.845 29.165 537.415 ;
  END
 END o317
 PIN o318
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 538.175 29.165 538.745 ;
  END
 END o318
 PIN o319
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 541.215 29.165 541.785 ;
  END
 END o319
 PIN o320
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 542.545 29.165 543.115 ;
  END
 END o320
 PIN o321
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 545.585 29.165 546.155 ;
  END
 END o321
 PIN o322
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 546.915 29.165 547.485 ;
  END
 END o322
 PIN o323
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 117.895 29.165 118.465 ;
  END
 END o323
 PIN o324
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 549.955 29.165 550.525 ;
  END
 END o324
 PIN o325
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 551.285 29.165 551.855 ;
  END
 END o325
 PIN o326
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 554.325 29.165 554.895 ;
  END
 END o326
 PIN o327
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 555.655 29.165 556.225 ;
  END
 END o327
 PIN o328
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 558.695 29.165 559.265 ;
  END
 END o328
 PIN o329
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 560.025 29.165 560.595 ;
  END
 END o329
 PIN o330
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 563.065 29.165 563.635 ;
  END
 END o330
 PIN o331
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 120.935 29.165 121.505 ;
  END
 END o331
 PIN o332
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 122.265 29.165 122.835 ;
  END
 END o332
 PIN o333
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 85.975 29.165 86.545 ;
  END
 END o333
 PIN o334
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 125.305 29.165 125.875 ;
  END
 END o334
 PIN o335
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 126.635 29.165 127.205 ;
  END
 END o335
 PIN o336
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 129.675 29.165 130.245 ;
  END
 END o336
 PIN o337
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 131.005 29.165 131.575 ;
  END
 END o337
 PIN o338
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 134.045 29.165 134.615 ;
  END
 END o338
 PIN o339
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 135.375 29.165 135.945 ;
  END
 END o339
 PIN o340
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 138.415 29.165 138.985 ;
  END
 END o340
 PIN o341
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 139.745 29.165 140.315 ;
  END
 END o341
 PIN o342
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 142.785 29.165 143.355 ;
  END
 END o342
 PIN o343
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 144.115 29.165 144.685 ;
  END
 END o343
 PIN o344
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 87.305 29.165 87.875 ;
  END
 END o344
 PIN o345
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 147.155 29.165 147.725 ;
  END
 END o345
 PIN o346
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 148.485 29.165 149.055 ;
  END
 END o346
 PIN o347
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 151.525 29.165 152.095 ;
  END
 END o347
 PIN o348
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 152.855 29.165 153.425 ;
  END
 END o348
 PIN o349
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 155.895 29.165 156.465 ;
  END
 END o349
 PIN o350
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 157.225 29.165 157.795 ;
  END
 END o350
 PIN o351
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 160.265 29.165 160.835 ;
  END
 END o351
 PIN o352
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 161.595 29.165 162.165 ;
  END
 END o352
 PIN o353
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 164.635 29.165 165.205 ;
  END
 END o353
 PIN o354
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 165.965 29.165 166.535 ;
  END
 END o354
 PIN o355
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 90.345 29.165 90.915 ;
  END
 END o355
 PIN o356
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 169.005 29.165 169.575 ;
  END
 END o356
 PIN o357
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 170.335 29.165 170.905 ;
  END
 END o357
 PIN o358
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 173.375 29.165 173.945 ;
  END
 END o358
 PIN o359
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 174.705 29.165 175.275 ;
  END
 END o359
 PIN o360
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 177.745 29.165 178.315 ;
  END
 END o360
 PIN o361
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 179.075 29.165 179.645 ;
  END
 END o361
 PIN o362
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 182.115 29.165 182.685 ;
  END
 END o362
 PIN o363
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 183.445 29.165 184.015 ;
  END
 END o363
 PIN o364
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 186.485 29.165 187.055 ;
  END
 END o364
 PIN o365
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 187.815 29.165 188.385 ;
  END
 END o365
 PIN o366
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 91.675 29.165 92.245 ;
  END
 END o366
 PIN o367
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 190.855 29.165 191.425 ;
  END
 END o367
 PIN o368
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 192.185 29.165 192.755 ;
  END
 END o368
 PIN o369
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 195.225 29.165 195.795 ;
  END
 END o369
 PIN o370
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 196.555 29.165 197.125 ;
  END
 END o370
 PIN o371
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 199.595 29.165 200.165 ;
  END
 END o371
 PIN o372
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 200.925 29.165 201.495 ;
  END
 END o372
 PIN o373
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 203.965 29.165 204.535 ;
  END
 END o373
 PIN o374
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 205.295 29.165 205.865 ;
  END
 END o374
 PIN o375
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 208.335 29.165 208.905 ;
  END
 END o375
 PIN o376
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 224.295 29.165 224.865 ;
  END
 END o376
 PIN o377
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 94.715 29.165 95.285 ;
  END
 END o377
 PIN o378
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 226.385 29.165 226.955 ;
  END
 END o378
 PIN o379
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 263.435 29.165 264.005 ;
  END
 END o379
 PIN o380
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 264.765 29.165 265.335 ;
  END
 END o380
 PIN o381
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 267.805 29.165 268.375 ;
  END
 END o381
 PIN o382
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 269.135 29.165 269.705 ;
  END
 END o382
 PIN o383
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 272.175 29.165 272.745 ;
  END
 END o383
 PIN o384
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 273.505 29.165 274.075 ;
  END
 END o384
 PIN o385
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 276.545 29.165 277.115 ;
  END
 END o385
 PIN o386
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 277.875 29.165 278.445 ;
  END
 END o386
 PIN o387
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 280.915 29.165 281.485 ;
  END
 END o387
 PIN o388
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 96.045 29.165 96.615 ;
  END
 END o388
 PIN o389
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 282.245 29.165 282.815 ;
  END
 END o389
 PIN o390
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 285.285 29.165 285.855 ;
  END
 END o390
 PIN o391
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 286.615 29.165 287.185 ;
  END
 END o391
 PIN o392
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 289.655 29.165 290.225 ;
  END
 END o392
 PIN o393
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 290.985 29.165 291.555 ;
  END
 END o393
 PIN o394
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 294.025 29.165 294.595 ;
  END
 END o394
 PIN o395
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 295.355 29.165 295.925 ;
  END
 END o395
 PIN o396
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 298.395 29.165 298.965 ;
  END
 END o396
 PIN o397
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 299.725 29.165 300.295 ;
  END
 END o397
 PIN o398
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 302.765 29.165 303.335 ;
  END
 END o398
 PIN o399
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 99.085 29.165 99.655 ;
  END
 END o399
 PIN o400
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 304.095 29.165 304.665 ;
  END
 END o400
 PIN o401
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 307.135 29.165 307.705 ;
  END
 END o401
 PIN o402
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 308.465 29.165 309.035 ;
  END
 END o402
 PIN o403
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 311.505 29.165 312.075 ;
  END
 END o403
 PIN o404
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 312.835 29.165 313.405 ;
  END
 END o404
 PIN o405
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 315.875 29.165 316.445 ;
  END
 END o405
 PIN o406
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 317.205 29.165 317.775 ;
  END
 END o406
 PIN o407
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 320.245 29.165 320.815 ;
  END
 END o407
 PIN o408
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 321.575 29.165 322.145 ;
  END
 END o408
 PIN o409
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 324.615 29.165 325.185 ;
  END
 END o409
 PIN o410
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 100.415 29.165 100.985 ;
  END
 END o410
 PIN o411
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 325.945 29.165 326.515 ;
  END
 END o411
 PIN o412
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 328.985 29.165 329.555 ;
  END
 END o412
 PIN o413
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 330.315 29.165 330.885 ;
  END
 END o413
 PIN o414
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 333.355 29.165 333.925 ;
  END
 END o414
 PIN o415
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 334.685 29.165 335.255 ;
  END
 END o415
 PIN o416
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 337.725 29.165 338.295 ;
  END
 END o416
 PIN o417
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 339.055 29.165 339.625 ;
  END
 END o417
 PIN o418
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 342.095 29.165 342.665 ;
  END
 END o418
 PIN o419
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 343.425 29.165 343.995 ;
  END
 END o419
 PIN o420
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 346.465 29.165 347.035 ;
  END
 END o420
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 54.815 0.665 55.385 1.235 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 44.175 0.665 44.745 1.235 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.575 0.665 56.145 1.235 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 42.275 0.665 42.845 1.235 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 56.335 0.665 56.905 1.235 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 43.415 0.665 43.985 1.235 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 345.895 10.925 346.465 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 341.525 10.925 342.095 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 339.435 10.925 340.005 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 337.155 10.925 337.725 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 49.115 10.925 49.685 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 553.945 10.925 554.515 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 551.665 10.925 552.235 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 549.575 10.925 550.145 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 352.545 10.925 353.115 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 350.265 10.925 350.835 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 348.175 10.925 348.745 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 343.805 10.925 344.375 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 332.785 10.925 333.355 ;
  END
 END i18
 PIN i19
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 328.415 10.925 328.985 ;
  END
 END i19
 PIN i20
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 321.955 10.925 322.525 ;
  END
 END i20
 PIN i21
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 335.065 10.925 335.635 ;
  END
 END i21
 PIN i22
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 326.325 10.925 326.895 ;
  END
 END i22
 PIN i23
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 98.705 10.925 99.275 ;
  END
 END i23
 PIN i24
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 313.215 10.925 313.785 ;
  END
 END i24
 PIN i25
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 310.935 10.925 311.505 ;
  END
 END i25
 PIN i26
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 308.845 10.925 309.415 ;
  END
 END i26
 PIN i27
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 306.565 10.925 307.135 ;
  END
 END i27
 PIN i28
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 302.195 10.925 302.765 ;
  END
 END i28
 PIN i29
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 300.105 10.925 300.675 ;
  END
 END i29
 PIN i30
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 297.825 10.925 298.395 ;
  END
 END i30
 PIN i31
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 96.425 10.925 96.995 ;
  END
 END i31
 PIN i32
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 304.475 10.925 305.045 ;
  END
 END i32
 PIN i33
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 100.795 10.925 101.365 ;
  END
 END i33
 PIN i34
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 319.675 10.925 320.245 ;
  END
 END i34
 PIN i35
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 317.585 10.925 318.155 ;
  END
 END i35
 PIN i36
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 315.305 10.925 315.875 ;
  END
 END i36
 PIN i37
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 135.755 10.925 136.325 ;
  END
 END i37
 PIN i38
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 129.295 10.925 129.865 ;
  END
 END i38
 PIN i39
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 131.385 10.925 131.955 ;
  END
 END i39
 PIN i40
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 133.665 10.925 134.235 ;
  END
 END i40
 PIN i41
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 124.925 10.925 125.495 ;
  END
 END i41
 PIN i42
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 127.015 10.925 127.585 ;
  END
 END i42
 PIN i43
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 122.645 10.925 123.215 ;
  END
 END i43
 PIN i44
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 47.025 10.925 47.595 ;
  END
 END i44
 PIN i45
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 89.965 10.925 90.535 ;
  END
 END i45
 PIN i46
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 545.205 10.925 545.775 ;
  END
 END i46
 PIN i47
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 547.295 10.925 547.865 ;
  END
 END i47
 PIN i48
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 111.815 10.925 112.385 ;
  END
 END i48
 PIN i49
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 523.355 10.925 523.925 ;
  END
 END i49
 PIN i50
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 512.335 10.925 512.905 ;
  END
 END i50
 PIN i51
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 113.905 10.925 114.475 ;
  END
 END i51
 PIN i52
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 148.865 10.925 149.435 ;
  END
 END i52
 PIN i53
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 116.185 10.925 116.755 ;
  END
 END i53
 PIN i54
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 120.555 10.925 121.125 ;
  END
 END i54
 PIN i55
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 374.395 10.925 374.965 ;
  END
 END i55
 PIN i56
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 118.275 10.925 118.845 ;
  END
 END i56
 PIN i57
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 85.595 10.925 86.165 ;
  END
 END i57
 PIN i58
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 138.035 10.925 138.605 ;
  END
 END i58
 PIN i59
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 361.285 10.925 361.855 ;
  END
 END i59
 PIN i60
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 383.135 10.925 383.705 ;
  END
 END i60
 PIN i61
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 363.375 10.925 363.945 ;
  END
 END i61
 PIN i62
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 560.405 10.925 560.975 ;
  END
 END i62
 PIN i63
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 558.315 10.925 558.885 ;
  END
 END i63
 PIN i64
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 403.845 10.925 404.415 ;
  END
 END i64
 PIN i65
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 359.005 10.925 359.575 ;
  END
 END i65
 PIN i66
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 401.755 10.925 402.325 ;
  END
 END i66
 PIN i67
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 556.035 10.925 556.605 ;
  END
 END i67
 PIN i68
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 380.855 10.925 381.425 ;
  END
 END i68
 PIN i69
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 103.075 10.925 103.645 ;
  END
 END i69
 PIN i70
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 365.655 10.925 366.225 ;
  END
 END i70
 PIN i71
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 105.165 10.925 105.735 ;
  END
 END i71
 PIN i72
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 109.535 10.925 110.105 ;
  END
 END i72
 PIN i73
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 354.635 10.925 355.205 ;
  END
 END i73
 PIN i74
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 295.735 10.925 296.305 ;
  END
 END i74
 PIN i75
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 177.365 10.925 177.935 ;
  END
 END i75
 PIN i76
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 510.245 10.925 510.815 ;
  END
 END i76
 PIN i77
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 501.505 10.925 502.075 ;
  END
 END i77
 PIN i78
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 521.075 10.925 521.645 ;
  END
 END i78
 PIN i79
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 516.705 10.925 517.275 ;
  END
 END i79
 PIN i80
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 518.985 10.925 519.555 ;
  END
 END i80
 PIN i81
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 525.445 10.925 526.015 ;
  END
 END i81
 PIN i82
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 464.265 10.925 464.835 ;
  END
 END i82
 PIN i83
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 470.915 10.925 471.485 ;
  END
 END i83
 PIN i84
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 440.325 10.925 440.895 ;
  END
 END i84
 PIN i85
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 161.975 10.925 162.545 ;
  END
 END i85
 PIN i86
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 155.515 10.925 156.085 ;
  END
 END i86
 PIN i87
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 144.495 10.925 145.065 ;
  END
 END i87
 PIN i88
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 140.125 10.925 140.695 ;
  END
 END i88
 PIN i89
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 367.745 10.925 368.315 ;
  END
 END i89
 PIN i90
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 457.805 10.925 458.375 ;
  END
 END i90
 PIN i91
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 376.485 10.925 377.055 ;
  END
 END i91
 PIN i92
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 107.445 10.925 108.015 ;
  END
 END i92
 PIN i93
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 372.115 10.925 372.685 ;
  END
 END i93
 PIN i94
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 378.765 10.925 379.335 ;
  END
 END i94
 PIN i95
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 278.255 10.925 278.825 ;
  END
 END i95
 PIN i96
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 275.975 10.925 276.545 ;
  END
 END i96
 PIN i97
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 282.625 10.925 283.195 ;
  END
 END i97
 PIN i98
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 271.605 10.925 272.175 ;
  END
 END i98
 PIN i99
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 289.085 10.925 289.655 ;
  END
 END i99
 PIN i100
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 192.565 10.925 193.135 ;
  END
 END i100
 PIN i101
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 194.845 10.925 195.415 ;
  END
 END i101
 PIN i102
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 190.475 10.925 191.045 ;
  END
 END i102
 PIN i103
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 179.455 10.925 180.025 ;
  END
 END i103
 PIN i104
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 181.735 10.925 182.305 ;
  END
 END i104
 PIN i105
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 172.995 10.925 173.565 ;
  END
 END i105
 PIN i106
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 183.825 10.925 184.395 ;
  END
 END i106
 PIN i107
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 186.105 10.925 186.675 ;
  END
 END i107
 PIN i108
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 170.715 10.925 171.285 ;
  END
 END i108
 PIN i109
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 175.085 10.925 175.655 ;
  END
 END i109
 PIN i110
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 188.195 10.925 188.765 ;
  END
 END i110
 PIN i111
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 540.835 10.925 541.405 ;
  END
 END i111
 PIN i112
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 538.555 10.925 539.125 ;
  END
 END i112
 PIN i113
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 507.965 10.925 508.535 ;
  END
 END i113
 PIN i114
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 505.875 10.925 506.445 ;
  END
 END i114
 PIN i115
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 497.135 10.925 497.705 ;
  END
 END i115
 PIN i116
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 494.855 10.925 495.425 ;
  END
 END i116
 PIN i117
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 486.115 10.925 486.685 ;
  END
 END i117
 PIN i118
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 503.595 10.925 504.165 ;
  END
 END i118
 PIN i119
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 490.485 10.925 491.055 ;
  END
 END i119
 PIN i120
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 492.765 10.925 493.335 ;
  END
 END i120
 PIN i121
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 499.225 10.925 499.795 ;
  END
 END i121
 PIN i122
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 488.395 10.925 488.965 ;
  END
 END i122
 PIN i123
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 536.465 10.925 537.035 ;
  END
 END i123
 PIN i124
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 534.185 10.925 534.755 ;
  END
 END i124
 PIN i125
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 527.725 10.925 528.295 ;
  END
 END i125
 PIN i126
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 514.615 10.925 515.185 ;
  END
 END i126
 PIN i127
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 532.095 10.925 532.665 ;
  END
 END i127
 PIN i128
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 459.895 10.925 460.465 ;
  END
 END i128
 PIN i129
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 462.175 10.925 462.745 ;
  END
 END i129
 PIN i130
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 466.545 10.925 467.115 ;
  END
 END i130
 PIN i131
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 468.635 10.925 469.205 ;
  END
 END i131
 PIN i132
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 455.525 10.925 456.095 ;
  END
 END i132
 PIN i133
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 151.145 10.925 151.715 ;
  END
 END i133
 PIN i134
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 442.415 10.925 442.985 ;
  END
 END i134
 PIN i135
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 451.155 10.925 451.725 ;
  END
 END i135
 PIN i136
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 475.285 10.925 475.855 ;
  END
 END i136
 PIN i137
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 481.745 10.925 482.315 ;
  END
 END i137
 PIN i138
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 446.785 10.925 447.355 ;
  END
 END i138
 PIN i139
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 484.025 10.925 484.595 ;
  END
 END i139
 PIN i140
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 153.235 10.925 153.805 ;
  END
 END i140
 PIN i141
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 479.655 10.925 480.225 ;
  END
 END i141
 PIN i142
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 157.605 10.925 158.175 ;
  END
 END i142
 PIN i143
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 164.255 10.925 164.825 ;
  END
 END i143
 PIN i144
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 473.005 10.925 473.575 ;
  END
 END i144
 PIN i145
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 453.435 10.925 454.005 ;
  END
 END i145
 PIN i146
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 542.925 10.925 543.495 ;
  END
 END i146
 PIN i147
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 529.815 10.925 530.385 ;
  END
 END i147
 PIN i148
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 477.375 10.925 477.945 ;
  END
 END i148
 PIN i149
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 356.915 10.925 357.485 ;
  END
 END i149
 PIN i150
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 87.685 10.925 88.255 ;
  END
 END i150
 PIN i151
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 203.585 10.925 204.155 ;
  END
 END i151
 PIN i152
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 205.675 10.925 206.245 ;
  END
 END i152
 PIN i153
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 166.345 10.925 166.915 ;
  END
 END i153
 PIN i154
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 207.955 10.925 208.525 ;
  END
 END i154
 PIN i155
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 226.575 10.925 227.145 ;
  END
 END i155
 PIN i156
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 280.345 10.925 280.915 ;
  END
 END i156
 PIN i157
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 286.995 10.925 287.565 ;
  END
 END i157
 PIN i158
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 146.775 10.925 147.345 ;
  END
 END i158
 PIN i159
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 262.865 10.925 263.435 ;
  END
 END i159
 PIN i160
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 267.235 10.925 267.805 ;
  END
 END i160
 PIN i161
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 269.515 10.925 270.085 ;
  END
 END i161
 PIN i162
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 291.365 10.925 291.935 ;
  END
 END i162
 PIN i163
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 92.055 10.925 92.625 ;
  END
 END i163
 PIN i164
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 94.335 10.925 94.905 ;
  END
 END i164
 PIN i165
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 142.405 10.925 142.975 ;
  END
 END i165
 PIN i166
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 168.625 10.925 169.195 ;
  END
 END i166
 PIN i167
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 196.935 10.925 197.505 ;
  END
 END i167
 PIN i168
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 199.215 10.925 199.785 ;
  END
 END i168
 PIN i169
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 201.305 10.925 201.875 ;
  END
 END i169
 PIN i170
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 224.295 10.925 224.865 ;
  END
 END i170
 PIN i171
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 265.145 10.925 265.715 ;
  END
 END i171
 PIN i172
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 273.885 10.925 274.455 ;
  END
 END i172
 PIN i173
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 284.715 10.925 285.285 ;
  END
 END i173
 PIN i174
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 293.455 10.925 294.025 ;
  END
 END i174
 PIN i175
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 324.045 10.925 324.615 ;
  END
 END i175
 PIN i176
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 330.695 10.925 331.265 ;
  END
 END i176
 PIN i177
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 370.025 10.925 370.595 ;
  END
 END i177
 PIN i178
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 449.065 10.925 449.635 ;
  END
 END i178
 PIN i179
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 159.885 10.925 160.455 ;
  END
 END i179
 PIN i180
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 444.695 10.925 445.265 ;
  END
 END i180
 PIN i181
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 385.225 10.925 385.795 ;
  END
 END i181
 PIN i182
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 59.375 0.665 59.945 1.235 ;
  END
 END i182
 PIN i183
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 37.715 0.665 38.285 1.235 ;
  END
 END i183
 PIN i184
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 35.815 0.665 36.385 1.235 ;
  END
 END i184
 PIN i185
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 60.895 0.665 61.465 1.235 ;
  END
 END i185
 PIN i186
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 39.615 0.665 40.185 1.235 ;
  END
 END i186
 PIN i187
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.295 0.665 34.865 1.235 ;
  END
 END i187
 PIN i188
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 70.015 0.665 70.585 1.235 ;
  END
 END i188
 PIN i189
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 0.665 71.725 1.235 ;
  END
 END i189
 PIN i190
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 38.855 0.665 39.425 1.235 ;
  END
 END i190
 PIN i191
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 62.035 0.665 62.605 1.235 ;
  END
 END i191
 PIN i192
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 60.135 0.665 60.705 1.235 ;
  END
 END i192
 PIN i193
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 35.055 0.665 35.625 1.235 ;
  END
 END i193
 PIN i194
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 36.955 0.665 37.525 1.235 ;
  END
 END i194
 PIN i195
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 47.025 4.085 47.595 ;
  END
 END i195
 PIN i196
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 48.735 4.085 49.305 ;
  END
 END i196
 PIN i197
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 103.265 4.085 103.835 ;
  END
 END i197
 PIN i198
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 347.795 4.085 348.365 ;
  END
 END i198
 PIN i199
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 350.455 4.085 351.025 ;
  END
 END i199
 PIN i200
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 352.165 4.085 352.735 ;
  END
 END i200
 PIN i201
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 354.825 4.085 355.395 ;
  END
 END i201
 PIN i202
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 356.535 4.085 357.105 ;
  END
 END i202
 PIN i203
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 359.195 4.085 359.765 ;
  END
 END i203
 PIN i204
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 360.905 4.085 361.475 ;
  END
 END i204
 PIN i205
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 363.565 4.085 364.135 ;
  END
 END i205
 PIN i206
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 365.275 4.085 365.845 ;
  END
 END i206
 PIN i207
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 367.935 4.085 368.505 ;
  END
 END i207
 PIN i208
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 104.975 4.085 105.545 ;
  END
 END i208
 PIN i209
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 369.645 4.085 370.215 ;
  END
 END i209
 PIN i210
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 372.305 4.085 372.875 ;
  END
 END i210
 PIN i211
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 374.015 4.085 374.585 ;
  END
 END i211
 PIN i212
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 376.675 4.085 377.245 ;
  END
 END i212
 PIN i213
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 378.385 4.085 378.955 ;
  END
 END i213
 PIN i214
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 381.045 4.085 381.615 ;
  END
 END i214
 PIN i215
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 382.755 4.085 383.325 ;
  END
 END i215
 PIN i216
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 385.415 4.085 385.985 ;
  END
 END i216
 PIN i217
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 401.565 4.085 402.135 ;
  END
 END i217
 PIN i218
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 403.275 4.085 403.845 ;
  END
 END i218
 PIN i219
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 107.635 4.085 108.205 ;
  END
 END i219
 PIN i220
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 440.515 4.085 441.085 ;
  END
 END i220
 PIN i221
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 442.225 4.085 442.795 ;
  END
 END i221
 PIN i222
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 444.885 4.085 445.455 ;
  END
 END i222
 PIN i223
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 446.595 4.085 447.165 ;
  END
 END i223
 PIN i224
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 449.255 4.085 449.825 ;
  END
 END i224
 PIN i225
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 450.965 4.085 451.535 ;
  END
 END i225
 PIN i226
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 453.625 4.085 454.195 ;
  END
 END i226
 PIN i227
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 455.335 4.085 455.905 ;
  END
 END i227
 PIN i228
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 457.995 4.085 458.565 ;
  END
 END i228
 PIN i229
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 459.705 4.085 460.275 ;
  END
 END i229
 PIN i230
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 109.345 4.085 109.915 ;
  END
 END i230
 PIN i231
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 462.365 4.085 462.935 ;
  END
 END i231
 PIN i232
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 464.075 4.085 464.645 ;
  END
 END i232
 PIN i233
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 466.735 4.085 467.305 ;
  END
 END i233
 PIN i234
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 468.445 4.085 469.015 ;
  END
 END i234
 PIN i235
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 471.105 4.085 471.675 ;
  END
 END i235
 PIN i236
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 472.815 4.085 473.385 ;
  END
 END i236
 PIN i237
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 475.475 4.085 476.045 ;
  END
 END i237
 PIN i238
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 477.185 4.085 477.755 ;
  END
 END i238
 PIN i239
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 479.845 4.085 480.415 ;
  END
 END i239
 PIN i240
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 481.555 4.085 482.125 ;
  END
 END i240
 PIN i241
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 112.005 4.085 112.575 ;
  END
 END i241
 PIN i242
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 484.215 4.085 484.785 ;
  END
 END i242
 PIN i243
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 485.925 4.085 486.495 ;
  END
 END i243
 PIN i244
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 488.585 4.085 489.155 ;
  END
 END i244
 PIN i245
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 490.295 4.085 490.865 ;
  END
 END i245
 PIN i246
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 492.955 4.085 493.525 ;
  END
 END i246
 PIN i247
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 494.665 4.085 495.235 ;
  END
 END i247
 PIN i248
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 497.325 4.085 497.895 ;
  END
 END i248
 PIN i249
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 499.035 4.085 499.605 ;
  END
 END i249
 PIN i250
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 501.695 4.085 502.265 ;
  END
 END i250
 PIN i251
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 503.405 4.085 503.975 ;
  END
 END i251
 PIN i252
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 113.715 4.085 114.285 ;
  END
 END i252
 PIN i253
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 506.065 4.085 506.635 ;
  END
 END i253
 PIN i254
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 507.775 4.085 508.345 ;
  END
 END i254
 PIN i255
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 510.435 4.085 511.005 ;
  END
 END i255
 PIN i256
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 512.145 4.085 512.715 ;
  END
 END i256
 PIN i257
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 514.805 4.085 515.375 ;
  END
 END i257
 PIN i258
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 516.515 4.085 517.085 ;
  END
 END i258
 PIN i259
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 519.175 4.085 519.745 ;
  END
 END i259
 PIN i260
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 520.885 4.085 521.455 ;
  END
 END i260
 PIN i261
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 523.545 4.085 524.115 ;
  END
 END i261
 PIN i262
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 525.255 4.085 525.825 ;
  END
 END i262
 PIN i263
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 116.375 4.085 116.945 ;
  END
 END i263
 PIN i264
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 527.915 4.085 528.485 ;
  END
 END i264
 PIN i265
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 529.625 4.085 530.195 ;
  END
 END i265
 PIN i266
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 532.285 4.085 532.855 ;
  END
 END i266
 PIN i267
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 533.995 4.085 534.565 ;
  END
 END i267
 PIN i268
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 536.655 4.085 537.225 ;
  END
 END i268
 PIN i269
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 538.365 4.085 538.935 ;
  END
 END i269
 PIN i270
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 541.025 4.085 541.595 ;
  END
 END i270
 PIN i271
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 542.735 4.085 543.305 ;
  END
 END i271
 PIN i272
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 545.395 4.085 545.965 ;
  END
 END i272
 PIN i273
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 547.105 4.085 547.675 ;
  END
 END i273
 PIN i274
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 118.085 4.085 118.655 ;
  END
 END i274
 PIN i275
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 549.765 4.085 550.335 ;
  END
 END i275
 PIN i276
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 551.475 4.085 552.045 ;
  END
 END i276
 PIN i277
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 554.135 4.085 554.705 ;
  END
 END i277
 PIN i278
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 555.845 4.085 556.415 ;
  END
 END i278
 PIN i279
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 558.505 4.085 559.075 ;
  END
 END i279
 PIN i280
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 560.215 4.085 560.785 ;
  END
 END i280
 PIN i281
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 562.875 4.085 563.445 ;
  END
 END i281
 PIN i282
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 120.745 4.085 121.315 ;
  END
 END i282
 PIN i283
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 122.455 4.085 123.025 ;
  END
 END i283
 PIN i284
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 85.785 4.085 86.355 ;
  END
 END i284
 PIN i285
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 125.115 4.085 125.685 ;
  END
 END i285
 PIN i286
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 126.825 4.085 127.395 ;
  END
 END i286
 PIN i287
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 129.485 4.085 130.055 ;
  END
 END i287
 PIN i288
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 131.195 4.085 131.765 ;
  END
 END i288
 PIN i289
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 133.855 4.085 134.425 ;
  END
 END i289
 PIN i290
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 135.565 4.085 136.135 ;
  END
 END i290
 PIN i291
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 138.225 4.085 138.795 ;
  END
 END i291
 PIN i292
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 139.935 4.085 140.505 ;
  END
 END i292
 PIN i293
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 142.595 4.085 143.165 ;
  END
 END i293
 PIN i294
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 144.305 4.085 144.875 ;
  END
 END i294
 PIN i295
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 87.495 4.085 88.065 ;
  END
 END i295
 PIN i296
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 146.965 4.085 147.535 ;
  END
 END i296
 PIN i297
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 148.675 4.085 149.245 ;
  END
 END i297
 PIN i298
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 151.335 4.085 151.905 ;
  END
 END i298
 PIN i299
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 153.045 4.085 153.615 ;
  END
 END i299
 PIN i300
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 155.705 4.085 156.275 ;
  END
 END i300
 PIN i301
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 157.415 4.085 157.985 ;
  END
 END i301
 PIN i302
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 160.075 4.085 160.645 ;
  END
 END i302
 PIN i303
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 161.785 4.085 162.355 ;
  END
 END i303
 PIN i304
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 164.445 4.085 165.015 ;
  END
 END i304
 PIN i305
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 166.155 4.085 166.725 ;
  END
 END i305
 PIN i306
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 90.155 4.085 90.725 ;
  END
 END i306
 PIN i307
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 168.815 4.085 169.385 ;
  END
 END i307
 PIN i308
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 170.525 4.085 171.095 ;
  END
 END i308
 PIN i309
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 173.185 4.085 173.755 ;
  END
 END i309
 PIN i310
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 174.895 4.085 175.465 ;
  END
 END i310
 PIN i311
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 177.555 4.085 178.125 ;
  END
 END i311
 PIN i312
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 179.265 4.085 179.835 ;
  END
 END i312
 PIN i313
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 181.925 4.085 182.495 ;
  END
 END i313
 PIN i314
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 183.635 4.085 184.205 ;
  END
 END i314
 PIN i315
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 186.295 4.085 186.865 ;
  END
 END i315
 PIN i316
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 188.005 4.085 188.575 ;
  END
 END i316
 PIN i317
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 91.865 4.085 92.435 ;
  END
 END i317
 PIN i318
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 190.665 4.085 191.235 ;
  END
 END i318
 PIN i319
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 192.375 4.085 192.945 ;
  END
 END i319
 PIN i320
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 195.035 4.085 195.605 ;
  END
 END i320
 PIN i321
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 196.745 4.085 197.315 ;
  END
 END i321
 PIN i322
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 199.405 4.085 199.975 ;
  END
 END i322
 PIN i323
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 201.115 4.085 201.685 ;
  END
 END i323
 PIN i324
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 203.775 4.085 204.345 ;
  END
 END i324
 PIN i325
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 205.485 4.085 206.055 ;
  END
 END i325
 PIN i326
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 208.145 4.085 208.715 ;
  END
 END i326
 PIN i327
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 224.295 4.085 224.865 ;
  END
 END i327
 PIN i328
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 94.525 4.085 95.095 ;
  END
 END i328
 PIN i329
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 226.005 4.085 226.575 ;
  END
 END i329
 PIN i330
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 263.055 4.085 263.625 ;
  END
 END i330
 PIN i331
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 264.765 4.085 265.335 ;
  END
 END i331
 PIN i332
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 267.425 4.085 267.995 ;
  END
 END i332
 PIN i333
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 269.135 4.085 269.705 ;
  END
 END i333
 PIN i334
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 271.795 4.085 272.365 ;
  END
 END i334
 PIN i335
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 273.505 4.085 274.075 ;
  END
 END i335
 PIN i336
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 276.165 4.085 276.735 ;
  END
 END i336
 PIN i337
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 277.875 4.085 278.445 ;
  END
 END i337
 PIN i338
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 280.535 4.085 281.105 ;
  END
 END i338
 PIN i339
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 96.235 4.085 96.805 ;
  END
 END i339
 PIN i340
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 282.245 4.085 282.815 ;
  END
 END i340
 PIN i341
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 284.905 4.085 285.475 ;
  END
 END i341
 PIN i342
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 286.615 4.085 287.185 ;
  END
 END i342
 PIN i343
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 289.275 4.085 289.845 ;
  END
 END i343
 PIN i344
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 290.985 4.085 291.555 ;
  END
 END i344
 PIN i345
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 293.645 4.085 294.215 ;
  END
 END i345
 PIN i346
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 295.355 4.085 295.925 ;
  END
 END i346
 PIN i347
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 298.015 4.085 298.585 ;
  END
 END i347
 PIN i348
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 299.725 4.085 300.295 ;
  END
 END i348
 PIN i349
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 302.385 4.085 302.955 ;
  END
 END i349
 PIN i350
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 98.895 4.085 99.465 ;
  END
 END i350
 PIN i351
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 304.095 4.085 304.665 ;
  END
 END i351
 PIN i352
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 306.755 4.085 307.325 ;
  END
 END i352
 PIN i353
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 308.465 4.085 309.035 ;
  END
 END i353
 PIN i354
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 311.125 4.085 311.695 ;
  END
 END i354
 PIN i355
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 312.835 4.085 313.405 ;
  END
 END i355
 PIN i356
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 315.495 4.085 316.065 ;
  END
 END i356
 PIN i357
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 317.205 4.085 317.775 ;
  END
 END i357
 PIN i358
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 319.865 4.085 320.435 ;
  END
 END i358
 PIN i359
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 321.575 4.085 322.145 ;
  END
 END i359
 PIN i360
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 324.235 4.085 324.805 ;
  END
 END i360
 PIN i361
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 100.605 4.085 101.175 ;
  END
 END i361
 PIN i362
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 325.945 4.085 326.515 ;
  END
 END i362
 PIN i363
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 328.605 4.085 329.175 ;
  END
 END i363
 PIN i364
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 330.315 4.085 330.885 ;
  END
 END i364
 PIN i365
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 332.975 4.085 333.545 ;
  END
 END i365
 PIN i366
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 334.685 4.085 335.255 ;
  END
 END i366
 PIN i367
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 337.345 4.085 337.915 ;
  END
 END i367
 PIN i368
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 339.055 4.085 339.625 ;
  END
 END i368
 PIN i369
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 341.715 4.085 342.285 ;
  END
 END i369
 PIN i370
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 343.425 4.085 343.995 ;
  END
 END i370
 PIN i371
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 346.085 4.085 346.655 ;
  END
 END i371
 PIN i372
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 46.455 3.325 47.025 ;
  END
 END i372
 PIN i373
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 49.115 3.325 49.685 ;
  END
 END i373
 PIN i374
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 102.695 3.325 103.265 ;
  END
 END i374
 PIN i375
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 348.365 3.325 348.935 ;
  END
 END i375
 PIN i376
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 350.075 3.325 350.645 ;
  END
 END i376
 PIN i377
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 352.735 3.325 353.305 ;
  END
 END i377
 PIN i378
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 354.445 3.325 355.015 ;
  END
 END i378
 PIN i379
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 357.105 3.325 357.675 ;
  END
 END i379
 PIN i380
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 358.815 3.325 359.385 ;
  END
 END i380
 PIN i381
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 361.475 3.325 362.045 ;
  END
 END i381
 PIN i382
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 363.185 3.325 363.755 ;
  END
 END i382
 PIN i383
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 365.845 3.325 366.415 ;
  END
 END i383
 PIN i384
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 367.555 3.325 368.125 ;
  END
 END i384
 PIN i385
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 105.355 3.325 105.925 ;
  END
 END i385
 PIN i386
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 370.215 3.325 370.785 ;
  END
 END i386
 PIN i387
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 371.925 3.325 372.495 ;
  END
 END i387
 PIN i388
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 374.585 3.325 375.155 ;
  END
 END i388
 PIN i389
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 376.295 3.325 376.865 ;
  END
 END i389
 PIN i390
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 378.955 3.325 379.525 ;
  END
 END i390
 PIN i391
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 380.665 3.325 381.235 ;
  END
 END i391
 PIN i392
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 383.325 3.325 383.895 ;
  END
 END i392
 PIN i393
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 385.035 3.325 385.605 ;
  END
 END i393
 PIN i394
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 401.185 3.325 401.755 ;
  END
 END i394
 PIN i395
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 403.845 3.325 404.415 ;
  END
 END i395
 PIN i396
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 107.065 3.325 107.635 ;
  END
 END i396
 PIN i397
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 439.945 3.325 440.515 ;
  END
 END i397
 PIN i398
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 442.605 3.325 443.175 ;
  END
 END i398
 PIN i399
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 444.315 3.325 444.885 ;
  END
 END i399
 PIN i400
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 446.975 3.325 447.545 ;
  END
 END i400
 PIN i401
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 448.685 3.325 449.255 ;
  END
 END i401
 PIN i402
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 451.345 3.325 451.915 ;
  END
 END i402
 PIN i403
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 453.055 3.325 453.625 ;
  END
 END i403
 PIN i404
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 455.715 3.325 456.285 ;
  END
 END i404
 PIN i405
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 457.425 3.325 457.995 ;
  END
 END i405
 PIN i406
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 460.085 3.325 460.655 ;
  END
 END i406
 PIN i407
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 109.725 3.325 110.295 ;
  END
 END i407
 PIN i408
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 461.795 3.325 462.365 ;
  END
 END i408
 PIN i409
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 464.455 3.325 465.025 ;
  END
 END i409
 PIN i410
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 466.165 3.325 466.735 ;
  END
 END i410
 PIN i411
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 468.825 3.325 469.395 ;
  END
 END i411
 PIN i412
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 470.535 3.325 471.105 ;
  END
 END i412
 PIN i413
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 473.195 3.325 473.765 ;
  END
 END i413
 PIN i414
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 474.905 3.325 475.475 ;
  END
 END i414
 PIN i415
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 477.565 3.325 478.135 ;
  END
 END i415
 PIN i416
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 479.275 3.325 479.845 ;
  END
 END i416
 PIN i417
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 481.935 3.325 482.505 ;
  END
 END i417
 PIN i418
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 111.435 3.325 112.005 ;
  END
 END i418
 PIN i419
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 483.645 3.325 484.215 ;
  END
 END i419
 PIN i420
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 486.305 3.325 486.875 ;
  END
 END i420
 PIN i421
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 488.015 3.325 488.585 ;
  END
 END i421
 PIN i422
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 490.675 3.325 491.245 ;
  END
 END i422
 PIN i423
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 492.385 3.325 492.955 ;
  END
 END i423
 PIN i424
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 495.045 3.325 495.615 ;
  END
 END i424
 PIN i425
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 496.755 3.325 497.325 ;
  END
 END i425
 PIN i426
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 499.415 3.325 499.985 ;
  END
 END i426
 PIN i427
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 501.125 3.325 501.695 ;
  END
 END i427
 PIN i428
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 503.785 3.325 504.355 ;
  END
 END i428
 PIN i429
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 114.095 3.325 114.665 ;
  END
 END i429
 PIN i430
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 505.495 3.325 506.065 ;
  END
 END i430
 PIN i431
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 508.155 3.325 508.725 ;
  END
 END i431
 PIN i432
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 509.865 3.325 510.435 ;
  END
 END i432
 PIN i433
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 512.525 3.325 513.095 ;
  END
 END i433
 PIN i434
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 514.235 3.325 514.805 ;
  END
 END i434
 PIN i435
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 516.895 3.325 517.465 ;
  END
 END i435
 PIN i436
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 518.605 3.325 519.175 ;
  END
 END i436
 PIN i437
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 521.265 3.325 521.835 ;
  END
 END i437
 PIN i438
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 522.975 3.325 523.545 ;
  END
 END i438
 PIN i439
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 525.635 3.325 526.205 ;
  END
 END i439
 PIN i440
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 115.805 3.325 116.375 ;
  END
 END i440
 PIN i441
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 527.345 3.325 527.915 ;
  END
 END i441
 PIN i442
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 530.005 3.325 530.575 ;
  END
 END i442
 PIN i443
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 531.715 3.325 532.285 ;
  END
 END i443
 PIN i444
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 534.375 3.325 534.945 ;
  END
 END i444
 PIN i445
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 536.085 3.325 536.655 ;
  END
 END i445
 PIN i446
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 538.745 3.325 539.315 ;
  END
 END i446
 PIN i447
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 540.455 3.325 541.025 ;
  END
 END i447
 PIN i448
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 543.115 3.325 543.685 ;
  END
 END i448
 PIN i449
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 544.825 3.325 545.395 ;
  END
 END i449
 PIN i450
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 547.485 3.325 548.055 ;
  END
 END i450
 PIN i451
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 118.465 3.325 119.035 ;
  END
 END i451
 PIN i452
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 549.195 3.325 549.765 ;
  END
 END i452
 PIN i453
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 551.855 3.325 552.425 ;
  END
 END i453
 PIN i454
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 553.565 3.325 554.135 ;
  END
 END i454
 PIN i455
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 556.225 3.325 556.795 ;
  END
 END i455
 PIN i456
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 557.935 3.325 558.505 ;
  END
 END i456
 PIN i457
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 560.595 3.325 561.165 ;
  END
 END i457
 PIN i458
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 562.305 3.325 562.875 ;
  END
 END i458
 PIN i459
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 120.175 3.325 120.745 ;
  END
 END i459
 PIN i460
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 122.835 3.325 123.405 ;
  END
 END i460
 PIN i461
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 85.215 3.325 85.785 ;
  END
 END i461
 PIN i462
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 124.545 3.325 125.115 ;
  END
 END i462
 PIN i463
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 127.205 3.325 127.775 ;
  END
 END i463
 PIN i464
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 128.915 3.325 129.485 ;
  END
 END i464
 PIN i465
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 131.575 3.325 132.145 ;
  END
 END i465
 PIN i466
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 133.285 3.325 133.855 ;
  END
 END i466
 PIN i467
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 135.945 3.325 136.515 ;
  END
 END i467
 PIN i468
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 137.655 3.325 138.225 ;
  END
 END i468
 PIN i469
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 140.315 3.325 140.885 ;
  END
 END i469
 PIN i470
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 142.025 3.325 142.595 ;
  END
 END i470
 PIN i471
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 144.685 3.325 145.255 ;
  END
 END i471
 PIN i472
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 87.875 3.325 88.445 ;
  END
 END i472
 PIN i473
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 146.395 3.325 146.965 ;
  END
 END i473
 PIN i474
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 149.055 3.325 149.625 ;
  END
 END i474
 PIN i475
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 150.765 3.325 151.335 ;
  END
 END i475
 PIN i476
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 153.425 3.325 153.995 ;
  END
 END i476
 PIN i477
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 155.135 3.325 155.705 ;
  END
 END i477
 PIN i478
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 157.795 3.325 158.365 ;
  END
 END i478
 PIN i479
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 159.505 3.325 160.075 ;
  END
 END i479
 PIN i480
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 162.165 3.325 162.735 ;
  END
 END i480
 PIN i481
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 163.875 3.325 164.445 ;
  END
 END i481
 PIN i482
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 166.535 3.325 167.105 ;
  END
 END i482
 PIN i483
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 89.585 3.325 90.155 ;
  END
 END i483
 PIN i484
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 168.245 3.325 168.815 ;
  END
 END i484
 PIN i485
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 170.905 3.325 171.475 ;
  END
 END i485
 PIN i486
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 172.615 3.325 173.185 ;
  END
 END i486
 PIN i487
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 175.275 3.325 175.845 ;
  END
 END i487
 PIN i488
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 176.985 3.325 177.555 ;
  END
 END i488
 PIN i489
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 179.645 3.325 180.215 ;
  END
 END i489
 PIN i490
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 181.355 3.325 181.925 ;
  END
 END i490
 PIN i491
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 184.015 3.325 184.585 ;
  END
 END i491
 PIN i492
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 185.725 3.325 186.295 ;
  END
 END i492
 PIN i493
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 188.385 3.325 188.955 ;
  END
 END i493
 PIN i494
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 92.245 3.325 92.815 ;
  END
 END i494
 PIN i495
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 190.095 3.325 190.665 ;
  END
 END i495
 PIN i496
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 192.755 3.325 193.325 ;
  END
 END i496
 PIN i497
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 194.465 3.325 195.035 ;
  END
 END i497
 PIN i498
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 197.125 3.325 197.695 ;
  END
 END i498
 PIN i499
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 198.835 3.325 199.405 ;
  END
 END i499
 PIN i500
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 201.495 3.325 202.065 ;
  END
 END i500
 PIN i501
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 203.205 3.325 203.775 ;
  END
 END i501
 PIN i502
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 205.865 3.325 206.435 ;
  END
 END i502
 PIN i503
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 207.575 3.325 208.145 ;
  END
 END i503
 PIN i504
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 223.725 3.325 224.295 ;
  END
 END i504
 PIN i505
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 93.955 3.325 94.525 ;
  END
 END i505
 PIN i506
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 226.385 3.325 226.955 ;
  END
 END i506
 PIN i507
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 262.675 3.325 263.245 ;
  END
 END i507
 PIN i508
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 265.335 3.325 265.905 ;
  END
 END i508
 PIN i509
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 267.045 3.325 267.615 ;
  END
 END i509
 PIN i510
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 269.705 3.325 270.275 ;
  END
 END i510
 PIN i511
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 271.415 3.325 271.985 ;
  END
 END i511
 PIN i512
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 274.075 3.325 274.645 ;
  END
 END i512
 PIN i513
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 275.785 3.325 276.355 ;
  END
 END i513
 PIN i514
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 278.445 3.325 279.015 ;
  END
 END i514
 PIN i515
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 280.155 3.325 280.725 ;
  END
 END i515
 PIN i516
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 96.615 3.325 97.185 ;
  END
 END i516
 PIN i517
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 282.815 3.325 283.385 ;
  END
 END i517
 PIN i518
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 284.525 3.325 285.095 ;
  END
 END i518
 PIN i519
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 287.185 3.325 287.755 ;
  END
 END i519
 PIN i520
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 288.895 3.325 289.465 ;
  END
 END i520
 PIN i521
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 291.555 3.325 292.125 ;
  END
 END i521
 PIN i522
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 293.265 3.325 293.835 ;
  END
 END i522
 PIN i523
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 295.925 3.325 296.495 ;
  END
 END i523
 PIN i524
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 297.635 3.325 298.205 ;
  END
 END i524
 PIN i525
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 300.295 3.325 300.865 ;
  END
 END i525
 PIN i526
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 302.005 3.325 302.575 ;
  END
 END i526
 PIN i527
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 98.325 3.325 98.895 ;
  END
 END i527
 PIN i528
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 304.665 3.325 305.235 ;
  END
 END i528
 PIN i529
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 306.375 3.325 306.945 ;
  END
 END i529
 PIN i530
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 309.035 3.325 309.605 ;
  END
 END i530
 PIN i531
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 310.745 3.325 311.315 ;
  END
 END i531
 PIN i532
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 313.405 3.325 313.975 ;
  END
 END i532
 PIN i533
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 315.115 3.325 315.685 ;
  END
 END i533
 PIN i534
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 317.775 3.325 318.345 ;
  END
 END i534
 PIN i535
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 319.485 3.325 320.055 ;
  END
 END i535
 PIN i536
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 322.145 3.325 322.715 ;
  END
 END i536
 PIN i537
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 323.855 3.325 324.425 ;
  END
 END i537
 PIN i538
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 100.985 3.325 101.555 ;
  END
 END i538
 PIN i539
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 326.515 3.325 327.085 ;
  END
 END i539
 PIN i540
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 328.225 3.325 328.795 ;
  END
 END i540
 PIN i541
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 330.885 3.325 331.455 ;
  END
 END i541
 PIN i542
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 332.595 3.325 333.165 ;
  END
 END i542
 PIN i543
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 335.255 3.325 335.825 ;
  END
 END i543
 PIN i544
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 336.965 3.325 337.535 ;
  END
 END i544
 PIN i545
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 339.625 3.325 340.195 ;
  END
 END i545
 PIN i546
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 341.335 3.325 341.905 ;
  END
 END i546
 PIN i547
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 343.995 3.325 344.565 ;
  END
 END i547
 PIN i548
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 345.705 3.325 346.275 ;
  END
 END i548
 PIN i549
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 65.455 3.325 66.025 ;
  END
 END i549
 PIN i550
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 242.725 3.325 243.295 ;
  END
 END i550
 PIN i551
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 420.185 3.325 420.755 ;
  END
 END i551
 PIN i552
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 46.075 4.085 46.645 ;
  END
 END i552
 PIN i553
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 49.685 4.085 50.255 ;
  END
 END i553
 PIN i554
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 102.315 4.085 102.885 ;
  END
 END i554
 PIN i555
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 348.745 4.085 349.315 ;
  END
 END i555
 PIN i556
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 349.505 4.085 350.075 ;
  END
 END i556
 PIN i557
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 353.115 4.085 353.685 ;
  END
 END i557
 PIN i558
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 353.875 4.085 354.445 ;
  END
 END i558
 PIN i559
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 357.485 4.085 358.055 ;
  END
 END i559
 PIN i560
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 358.245 4.085 358.815 ;
  END
 END i560
 PIN i561
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 361.855 4.085 362.425 ;
  END
 END i561
 PIN i562
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 362.615 4.085 363.185 ;
  END
 END i562
 PIN i563
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 366.225 4.085 366.795 ;
  END
 END i563
 PIN i564
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 366.985 4.085 367.555 ;
  END
 END i564
 PIN i565
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 105.925 4.085 106.495 ;
  END
 END i565
 PIN i566
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 370.595 4.085 371.165 ;
  END
 END i566
 PIN i567
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 371.355 4.085 371.925 ;
  END
 END i567
 PIN i568
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 374.965 4.085 375.535 ;
  END
 END i568
 PIN i569
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 375.725 4.085 376.295 ;
  END
 END i569
 PIN i570
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 379.335 4.085 379.905 ;
  END
 END i570
 PIN i571
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 380.095 4.085 380.665 ;
  END
 END i571
 PIN i572
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 383.705 4.085 384.275 ;
  END
 END i572
 PIN i573
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 384.465 4.085 385.035 ;
  END
 END i573
 PIN i574
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 400.615 4.085 401.185 ;
  END
 END i574
 PIN i575
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 404.225 4.085 404.795 ;
  END
 END i575
 PIN i576
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 106.685 4.085 107.255 ;
  END
 END i576
 PIN i577
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 439.565 4.085 440.135 ;
  END
 END i577
 PIN i578
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 443.175 4.085 443.745 ;
  END
 END i578
 PIN i579
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 443.935 4.085 444.505 ;
  END
 END i579
 PIN i580
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 447.545 4.085 448.115 ;
  END
 END i580
 PIN i581
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 448.305 4.085 448.875 ;
  END
 END i581
 PIN i582
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 451.915 4.085 452.485 ;
  END
 END i582
 PIN i583
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 452.675 4.085 453.245 ;
  END
 END i583
 PIN i584
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 456.285 4.085 456.855 ;
  END
 END i584
 PIN i585
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 457.045 4.085 457.615 ;
  END
 END i585
 PIN i586
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 460.655 4.085 461.225 ;
  END
 END i586
 PIN i587
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 110.295 4.085 110.865 ;
  END
 END i587
 PIN i588
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 461.415 4.085 461.985 ;
  END
 END i588
 PIN i589
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 465.025 4.085 465.595 ;
  END
 END i589
 PIN i590
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 465.785 4.085 466.355 ;
  END
 END i590
 PIN i591
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 469.395 4.085 469.965 ;
  END
 END i591
 PIN i592
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 470.155 4.085 470.725 ;
  END
 END i592
 PIN i593
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 473.765 4.085 474.335 ;
  END
 END i593
 PIN i594
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 474.525 4.085 475.095 ;
  END
 END i594
 PIN i595
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 478.135 4.085 478.705 ;
  END
 END i595
 PIN i596
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 478.895 4.085 479.465 ;
  END
 END i596
 PIN i597
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 482.505 4.085 483.075 ;
  END
 END i597
 PIN i598
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 111.055 4.085 111.625 ;
  END
 END i598
 PIN i599
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 483.265 4.085 483.835 ;
  END
 END i599
 PIN i600
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 486.875 4.085 487.445 ;
  END
 END i600
 PIN i601
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 487.635 4.085 488.205 ;
  END
 END i601
 PIN i602
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 491.245 4.085 491.815 ;
  END
 END i602
 PIN i603
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 492.005 4.085 492.575 ;
  END
 END i603
 PIN i604
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 495.615 4.085 496.185 ;
  END
 END i604
 PIN i605
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 496.375 4.085 496.945 ;
  END
 END i605
 PIN i606
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 499.985 4.085 500.555 ;
  END
 END i606
 PIN i607
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 500.745 4.085 501.315 ;
  END
 END i607
 PIN i608
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 504.355 4.085 504.925 ;
  END
 END i608
 PIN i609
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 114.665 4.085 115.235 ;
  END
 END i609
 PIN i610
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 505.115 4.085 505.685 ;
  END
 END i610
 PIN i611
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 508.725 4.085 509.295 ;
  END
 END i611
 PIN i612
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 509.485 4.085 510.055 ;
  END
 END i612
 PIN i613
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 513.095 4.085 513.665 ;
  END
 END i613
 PIN i614
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 513.855 4.085 514.425 ;
  END
 END i614
 PIN i615
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 517.465 4.085 518.035 ;
  END
 END i615
 PIN i616
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 518.225 4.085 518.795 ;
  END
 END i616
 PIN i617
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 521.835 4.085 522.405 ;
  END
 END i617
 PIN i618
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 522.595 4.085 523.165 ;
  END
 END i618
 PIN i619
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 526.205 4.085 526.775 ;
  END
 END i619
 PIN i620
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 115.425 4.085 115.995 ;
  END
 END i620
 PIN i621
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 526.965 4.085 527.535 ;
  END
 END i621
 PIN i622
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 530.575 4.085 531.145 ;
  END
 END i622
 PIN i623
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 531.335 4.085 531.905 ;
  END
 END i623
 PIN i624
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 534.945 4.085 535.515 ;
  END
 END i624
 PIN i625
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 535.705 4.085 536.275 ;
  END
 END i625
 PIN i626
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 539.315 4.085 539.885 ;
  END
 END i626
 PIN i627
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 540.075 4.085 540.645 ;
  END
 END i627
 PIN i628
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 543.685 4.085 544.255 ;
  END
 END i628
 PIN i629
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 544.445 4.085 545.015 ;
  END
 END i629
 PIN i630
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 548.055 4.085 548.625 ;
  END
 END i630
 PIN i631
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 119.035 4.085 119.605 ;
  END
 END i631
 PIN i632
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 548.815 4.085 549.385 ;
  END
 END i632
 PIN i633
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 552.425 4.085 552.995 ;
  END
 END i633
 PIN i634
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 553.185 4.085 553.755 ;
  END
 END i634
 PIN i635
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 556.795 4.085 557.365 ;
  END
 END i635
 PIN i636
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 557.555 4.085 558.125 ;
  END
 END i636
 PIN i637
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 561.165 4.085 561.735 ;
  END
 END i637
 PIN i638
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 561.925 4.085 562.495 ;
  END
 END i638
 PIN i639
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 119.795 4.085 120.365 ;
  END
 END i639
 PIN i640
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 123.405 4.085 123.975 ;
  END
 END i640
 PIN i641
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 84.835 4.085 85.405 ;
  END
 END i641
 PIN i642
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 124.165 4.085 124.735 ;
  END
 END i642
 PIN i643
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 127.775 4.085 128.345 ;
  END
 END i643
 PIN i644
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 128.535 4.085 129.105 ;
  END
 END i644
 PIN i645
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 132.145 4.085 132.715 ;
  END
 END i645
 PIN i646
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 132.905 4.085 133.475 ;
  END
 END i646
 PIN i647
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 136.515 4.085 137.085 ;
  END
 END i647
 PIN i648
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 137.275 4.085 137.845 ;
  END
 END i648
 PIN i649
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 140.885 4.085 141.455 ;
  END
 END i649
 PIN i650
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 141.645 4.085 142.215 ;
  END
 END i650
 PIN i651
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 145.255 4.085 145.825 ;
  END
 END i651
 PIN i652
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 88.445 4.085 89.015 ;
  END
 END i652
 PIN i653
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 146.015 4.085 146.585 ;
  END
 END i653
 PIN i654
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 149.625 4.085 150.195 ;
  END
 END i654
 PIN i655
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 150.385 4.085 150.955 ;
  END
 END i655
 PIN i656
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 153.995 4.085 154.565 ;
  END
 END i656
 PIN i657
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 154.755 4.085 155.325 ;
  END
 END i657
 PIN i658
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 158.365 4.085 158.935 ;
  END
 END i658
 PIN i659
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 159.125 4.085 159.695 ;
  END
 END i659
 PIN i660
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 162.735 4.085 163.305 ;
  END
 END i660
 PIN i661
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 163.495 4.085 164.065 ;
  END
 END i661
 PIN i662
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 167.105 4.085 167.675 ;
  END
 END i662
 PIN i663
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 89.205 4.085 89.775 ;
  END
 END i663
 PIN i664
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 167.865 4.085 168.435 ;
  END
 END i664
 PIN i665
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 171.475 4.085 172.045 ;
  END
 END i665
 PIN i666
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 172.235 4.085 172.805 ;
  END
 END i666
 PIN i667
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 175.845 4.085 176.415 ;
  END
 END i667
 PIN i668
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 176.605 4.085 177.175 ;
  END
 END i668
 PIN i669
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 180.215 4.085 180.785 ;
  END
 END i669
 PIN i670
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 180.975 4.085 181.545 ;
  END
 END i670
 PIN i671
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 184.585 4.085 185.155 ;
  END
 END i671
 PIN i672
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 185.345 4.085 185.915 ;
  END
 END i672
 PIN i673
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 188.955 4.085 189.525 ;
  END
 END i673
 PIN i674
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 92.815 4.085 93.385 ;
  END
 END i674
 PIN i675
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 189.715 4.085 190.285 ;
  END
 END i675
 PIN i676
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 193.325 4.085 193.895 ;
  END
 END i676
 PIN i677
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 194.085 4.085 194.655 ;
  END
 END i677
 PIN i678
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 197.695 4.085 198.265 ;
  END
 END i678
 PIN i679
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 198.455 4.085 199.025 ;
  END
 END i679
 PIN i680
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 202.065 4.085 202.635 ;
  END
 END i680
 PIN i681
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 202.825 4.085 203.395 ;
  END
 END i681
 PIN i682
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 206.435 4.085 207.005 ;
  END
 END i682
 PIN i683
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 207.195 4.085 207.765 ;
  END
 END i683
 PIN i684
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 223.345 4.085 223.915 ;
  END
 END i684
 PIN i685
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 93.575 4.085 94.145 ;
  END
 END i685
 PIN i686
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 226.955 4.085 227.525 ;
  END
 END i686
 PIN i687
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 262.105 4.085 262.675 ;
  END
 END i687
 PIN i688
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 265.715 4.085 266.285 ;
  END
 END i688
 PIN i689
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 266.475 4.085 267.045 ;
  END
 END i689
 PIN i690
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 270.085 4.085 270.655 ;
  END
 END i690
 PIN i691
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 270.845 4.085 271.415 ;
  END
 END i691
 PIN i692
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 274.455 4.085 275.025 ;
  END
 END i692
 PIN i693
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 275.215 4.085 275.785 ;
  END
 END i693
 PIN i694
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 278.825 4.085 279.395 ;
  END
 END i694
 PIN i695
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 279.585 4.085 280.155 ;
  END
 END i695
 PIN i696
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 97.185 4.085 97.755 ;
  END
 END i696
 PIN i697
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 283.195 4.085 283.765 ;
  END
 END i697
 PIN i698
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 283.955 4.085 284.525 ;
  END
 END i698
 PIN i699
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 287.565 4.085 288.135 ;
  END
 END i699
 PIN i700
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 288.325 4.085 288.895 ;
  END
 END i700
 PIN i701
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 291.935 4.085 292.505 ;
  END
 END i701
 PIN i702
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 292.695 4.085 293.265 ;
  END
 END i702
 PIN i703
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 296.305 4.085 296.875 ;
  END
 END i703
 PIN i704
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 297.065 4.085 297.635 ;
  END
 END i704
 PIN i705
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 300.675 4.085 301.245 ;
  END
 END i705
 PIN i706
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 301.435 4.085 302.005 ;
  END
 END i706
 PIN i707
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 97.945 4.085 98.515 ;
  END
 END i707
 PIN i708
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 305.045 4.085 305.615 ;
  END
 END i708
 PIN i709
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 305.805 4.085 306.375 ;
  END
 END i709
 PIN i710
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 309.415 4.085 309.985 ;
  END
 END i710
 PIN i711
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 310.175 4.085 310.745 ;
  END
 END i711
 PIN i712
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 313.785 4.085 314.355 ;
  END
 END i712
 PIN i713
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 314.545 4.085 315.115 ;
  END
 END i713
 PIN i714
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 318.155 4.085 318.725 ;
  END
 END i714
 PIN i715
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 318.915 4.085 319.485 ;
  END
 END i715
 PIN i716
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 322.525 4.085 323.095 ;
  END
 END i716
 PIN i717
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 323.285 4.085 323.855 ;
  END
 END i717
 PIN i718
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 101.555 4.085 102.125 ;
  END
 END i718
 PIN i719
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 326.895 4.085 327.465 ;
  END
 END i719
 PIN i720
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 327.655 4.085 328.225 ;
  END
 END i720
 PIN i721
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 331.265 4.085 331.835 ;
  END
 END i721
 PIN i722
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 332.025 4.085 332.595 ;
  END
 END i722
 PIN i723
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 335.635 4.085 336.205 ;
  END
 END i723
 PIN i724
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 336.395 4.085 336.965 ;
  END
 END i724
 PIN i725
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 340.005 4.085 340.575 ;
  END
 END i725
 PIN i726
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 340.765 4.085 341.335 ;
  END
 END i726
 PIN i727
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 344.375 4.085 344.945 ;
  END
 END i727
 PIN i728
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 345.135 4.085 345.705 ;
  END
 END i728
 PIN i729
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 69.255 0.665 69.825 1.235 ;
  END
 END i729
 PIN i730
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 63.935 0.665 64.505 1.235 ;
  END
 END i730
 PIN i731
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 64.695 0.665 65.265 1.235 ;
  END
 END i731
 PIN i732
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 65.455 0.665 66.025 1.235 ;
  END
 END i732
 PIN i733
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 66.595 0.665 67.165 1.235 ;
  END
 END i733
 PIN i734
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 67.355 0.665 67.925 1.235 ;
  END
 END i734
 PIN i735
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 68.495 0.665 69.065 1.235 ;
  END
 END i735
 PIN i736
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 74.575 0.665 75.145 1.235 ;
  END
 END i736
 PIN i737
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 44.935 0.665 45.505 1.235 ;
  END
 END i737
 PIN i738
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 53.675 0.665 54.245 1.235 ;
  END
 END i738
 PIN i739
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 46.075 0.665 46.645 1.235 ;
  END
 END i739
 PIN i740
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 52.915 0.665 53.485 1.235 ;
  END
 END i740
 PIN i741
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 46.835 0.665 47.405 1.235 ;
  END
 END i741
 PIN i742
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 51.775 0.665 52.345 1.235 ;
  END
 END i742
 PIN i743
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 101.175 0.665 101.745 1.235 ;
  END
 END i743
 PIN i744
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 104.595 0.665 105.165 1.235 ;
  END
 END i744
 PIN i745
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 120.175 0.665 120.745 1.235 ;
  END
 END i745
 PIN i746
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 124.735 0.665 125.305 1.235 ;
  END
 END i746
 PIN i747
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 126.635 0.665 127.205 1.235 ;
  END
 END i747
 PIN i748
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.295 0.665 129.865 1.235 ;
  END
 END i748
 PIN i749
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 131.195 0.665 131.765 1.235 ;
  END
 END i749
 PIN i750
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 95.855 0.665 96.425 1.235 ;
  END
 END i750
 PIN i751
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 92.815 0.665 93.385 1.235 ;
  END
 END i751
 PIN i752
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 90.155 0.665 90.725 1.235 ;
  END
 END i752
 PIN i753
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 85.595 0.665 86.165 1.235 ;
  END
 END i753
 PIN i754
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 119.415 0.665 119.985 1.235 ;
  END
 END i754
 PIN i755
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 109.155 0.665 109.725 1.235 ;
  END
 END i755
 PIN i756
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 112.955 0.665 113.525 1.235 ;
  END
 END i756
 PIN i757
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 116.755 0.665 117.325 1.235 ;
  END
 END i757
 PIN i758
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 112.195 0.665 112.765 1.235 ;
  END
 END i758
 PIN i759
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 108.395 0.665 108.965 1.235 ;
  END
 END i759
 PIN i760
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 103.835 0.665 104.405 1.235 ;
  END
 END i760
 PIN i761
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 100.035 0.665 100.605 1.235 ;
  END
 END i761
 PIN i762
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 115.615 0.665 116.185 1.235 ;
  END
 END i762
 PIN i763
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 77.995 0.665 78.565 1.235 ;
  END
 END i763
 PIN i764
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 79.135 0.665 79.705 1.235 ;
  END
 END i764
 PIN i765
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 81.795 0.665 82.365 1.235 ;
  END
 END i765
 PIN i766
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 82.935 0.665 83.505 1.235 ;
  END
 END i766
 PIN i767
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 86.355 0.665 86.925 1.235 ;
  END
 END i767
 PIN i768
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 87.495 0.665 88.065 1.235 ;
  END
 END i768
 PIN i769
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 89.015 0.665 89.585 1.235 ;
  END
 END i769
 PIN i770
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 76.095 0.665 76.665 1.235 ;
  END
 END i770
 OBS
  LAYER metal1 ;
   RECT 0 0 280.06 584.82 ;
  LAYER via1 ;
   RECT 0 0 280.06 584.82 ;
  LAYER metal2 ;
   RECT 0 0 280.06 584.82 ;
  LAYER via2 ;
   RECT 0 0 280.06 584.82 ;
  LAYER metal3 ;
   RECT 0 0 280.06 584.82 ;
  LAYER via3 ;
   RECT 0 0 280.06 584.82 ;
  LAYER metal4 ;
   RECT 0 0 280.06 584.82 ;
 END
END block_737x3078_1192

MACRO block_644x675_93
 CLASS BLOCK ;
 FOREIGN block_644x675_93 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 244.72 BY 128.25 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 33.535 241.585 34.105 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 33.915 240.825 34.485 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 34.295 241.585 34.865 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 34.675 240.825 35.245 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 35.055 241.585 35.625 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 35.435 240.825 36.005 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 35.815 241.585 36.385 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 36.195 240.825 36.765 ;
  END
 END o7
 PIN o8
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 36.575 241.585 37.145 ;
  END
 END o8
 PIN o9
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 36.955 240.825 37.525 ;
  END
 END o9
 PIN o10
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 38.095 241.585 38.665 ;
  END
 END o10
 PIN o11
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 38.475 240.825 39.045 ;
  END
 END o11
 PIN o12
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 38.855 241.585 39.425 ;
  END
 END o12
 PIN o13
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 39.235 240.825 39.805 ;
  END
 END o13
 PIN o14
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 39.615 241.585 40.185 ;
  END
 END o14
 PIN o15
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 39.995 240.825 40.565 ;
  END
 END o15
 PIN o16
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 40.375 241.585 40.945 ;
  END
 END o16
 PIN o17
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 40.755 240.825 41.325 ;
  END
 END o17
 PIN o18
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 41.135 241.585 41.705 ;
  END
 END o18
 PIN o19
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 43.415 241.585 43.985 ;
  END
 END o19
 PIN o20
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 43.795 240.825 44.365 ;
  END
 END o20
 PIN o21
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 44.175 241.585 44.745 ;
  END
 END o21
 PIN o22
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 44.555 240.825 45.125 ;
  END
 END o22
 PIN o23
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 44.935 241.585 45.505 ;
  END
 END o23
 PIN o24
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 45.315 240.825 45.885 ;
  END
 END o24
 PIN o25
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 45.695 241.585 46.265 ;
  END
 END o25
 PIN o26
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 46.075 240.825 46.645 ;
  END
 END o26
 PIN o27
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 47.215 241.585 47.785 ;
  END
 END o27
 PIN o28
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 47.595 240.825 48.165 ;
  END
 END o28
 PIN o29
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 47.975 241.585 48.545 ;
  END
 END o29
 PIN o30
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 48.355 240.825 48.925 ;
  END
 END o30
 PIN o31
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 48.735 241.585 49.305 ;
  END
 END o31
 PIN o32
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 49.495 241.585 50.065 ;
  END
 END o32
 PIN o33
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 49.875 240.825 50.445 ;
  END
 END o33
 PIN o34
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 50.255 241.585 50.825 ;
  END
 END o34
 PIN o35
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 68.115 241.585 68.685 ;
  END
 END o35
 PIN o36
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 68.875 241.585 69.445 ;
  END
 END o36
 PIN o37
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 70.395 241.585 70.965 ;
  END
 END o37
 PIN o38
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 70.775 240.825 71.345 ;
  END
 END o38
 PIN o39
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 71.155 241.585 71.725 ;
  END
 END o39
 PIN o40
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 71.535 240.825 72.105 ;
  END
 END o40
 PIN o41
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 50.635 240.825 51.205 ;
  END
 END o41
 PIN o42
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 52.535 241.585 53.105 ;
  END
 END o42
 PIN o43
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 52.915 240.825 53.485 ;
  END
 END o43
 PIN o44
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 53.675 241.585 54.245 ;
  END
 END o44
 PIN o45
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 54.055 240.825 54.625 ;
  END
 END o45
 PIN o46
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 54.435 241.585 55.005 ;
  END
 END o46
 PIN o47
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 54.815 240.825 55.385 ;
  END
 END o47
 PIN o48
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 55.195 241.585 55.765 ;
  END
 END o48
 PIN o49
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 56.335 241.585 56.905 ;
  END
 END o49
 PIN o50
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 56.715 240.825 57.285 ;
  END
 END o50
 PIN o51
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 57.095 241.585 57.665 ;
  END
 END o51
 PIN o52
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 57.475 240.825 58.045 ;
  END
 END o52
 PIN o53
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 57.855 241.585 58.425 ;
  END
 END o53
 PIN o54
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 58.235 240.825 58.805 ;
  END
 END o54
 PIN o55
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 58.615 241.585 59.185 ;
  END
 END o55
 PIN o56
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 58.995 240.825 59.565 ;
  END
 END o56
 PIN o57
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 59.375 241.585 59.945 ;
  END
 END o57
 PIN o58
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 240.255 59.755 240.825 60.325 ;
  END
 END o58
 PIN o59
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 63.935 124.545 64.505 125.115 ;
  END
 END o59
 PIN o60
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 67.355 124.545 67.925 125.115 ;
  END
 END o60
 PIN o61
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 80.655 124.545 81.225 125.115 ;
  END
 END o61
 PIN o62
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 98.515 124.545 99.085 125.115 ;
  END
 END o62
 PIN o63
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 48.355 3.325 48.925 ;
  END
 END o63
 PIN o64
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 40.375 3.325 40.945 ;
  END
 END o64
 PIN o65
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 39.615 3.325 40.185 ;
  END
 END o65
 PIN o66
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 47.975 4.085 48.545 ;
  END
 END o66
 PIN o67
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 44.935 3.325 45.505 ;
  END
 END o67
 PIN o68
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 44.175 3.325 44.745 ;
  END
 END o68
 PIN o69
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.675 124.545 130.245 125.115 ;
  END
 END o69
 PIN o70
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 135.375 124.545 135.945 125.115 ;
  END
 END o70
 PIN o71
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 168.435 124.545 169.005 125.115 ;
  END
 END o71
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 37.335 124.545 37.905 125.115 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 33.915 124.545 34.485 125.115 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 36.195 124.545 36.765 125.115 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 43.795 124.545 44.365 125.115 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 51.775 124.545 52.345 125.115 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 52.915 124.545 53.485 125.115 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 54.815 124.545 55.385 125.115 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 56.335 124.545 56.905 125.115 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 57.475 124.545 58.045 125.115 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 59.375 124.545 59.945 125.115 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 60.515 124.545 61.085 125.115 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 47.215 124.545 47.785 125.115 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 49.495 124.545 50.065 125.115 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 48.355 124.545 48.925 125.115 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 65.075 124.545 65.645 125.115 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 96.235 124.545 96.805 125.115 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 127.395 124.545 127.965 125.115 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 166.155 124.545 166.725 125.115 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 60.895 241.585 61.465 ;
  END
 END i18
 PIN i19
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 63.935 241.585 64.505 ;
  END
 END i19
 PIN i20
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 63.935 3.325 64.505 ;
  END
 END i20
 OBS
  LAYER metal1 ;
   RECT 0 0 244.72 128.25 ;
  LAYER via1 ;
   RECT 0 0 244.72 128.25 ;
  LAYER metal2 ;
   RECT 0 0 244.72 128.25 ;
  LAYER via2 ;
   RECT 0 0 244.72 128.25 ;
  LAYER metal3 ;
   RECT 0 0 244.72 128.25 ;
  LAYER via3 ;
   RECT 0 0 244.72 128.25 ;
  LAYER metal4 ;
   RECT 0 0 244.72 128.25 ;
 END
END block_644x675_93

MACRO block_321x324_65
 CLASS BLOCK ;
 FOREIGN block_321x324_65 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 121.98 BY 61.56 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 44.175 118.845 44.745 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 34.295 3.325 34.865 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 35.815 3.325 36.385 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 38.095 3.325 38.665 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 39.615 3.325 40.185 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 41.135 3.325 41.705 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 42.655 3.325 43.225 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 44.175 3.325 44.745 ;
  END
 END o7
 PIN o8
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 45.695 3.325 46.265 ;
  END
 END o8
 PIN o9
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 22.895 118.845 23.465 ;
  END
 END o9
 PIN o10
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 6.935 3.325 7.505 ;
  END
 END o10
 PIN o11
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 7.695 3.325 8.265 ;
  END
 END o11
 PIN o12
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 19.855 3.325 20.425 ;
  END
 END o12
 PIN o13
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 21.375 3.325 21.945 ;
  END
 END o13
 PIN o14
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 22.135 3.325 22.705 ;
  END
 END o14
 PIN o15
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 24.415 3.325 24.985 ;
  END
 END o15
 PIN o16
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 25.935 3.325 26.505 ;
  END
 END o16
 PIN o17
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 26.695 3.325 27.265 ;
  END
 END o17
 PIN o18
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 27.455 3.325 28.025 ;
  END
 END o18
 PIN o19
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 28.975 3.325 29.545 ;
  END
 END o19
 PIN o20
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 30.495 3.325 31.065 ;
  END
 END o20
 PIN o21
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 32.015 3.325 32.585 ;
  END
 END o21
 PIN o22
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 9.215 3.325 9.785 ;
  END
 END o22
 PIN o23
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 10.735 3.325 11.305 ;
  END
 END o23
 PIN o24
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 11.495 3.325 12.065 ;
  END
 END o24
 PIN o25
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 12.255 3.325 12.825 ;
  END
 END o25
 PIN o26
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 13.775 3.325 14.345 ;
  END
 END o26
 PIN o27
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 15.295 3.325 15.865 ;
  END
 END o27
 PIN o28
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 16.055 3.325 16.625 ;
  END
 END o28
 PIN o29
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 16.815 3.325 17.385 ;
  END
 END o29
 PIN o30
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 25.175 118.845 25.745 ;
  END
 END o30
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 32.015 118.845 32.585 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 44.935 118.845 45.505 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 30.495 118.845 31.065 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 31.255 118.845 31.825 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 35.055 118.845 35.625 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 34.295 118.845 34.865 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 27.455 118.845 28.025 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 28.975 118.845 29.545 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 24.415 118.845 24.985 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 42.655 118.845 43.225 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 47.215 3.325 47.785 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 4.655 3.325 5.225 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 22.135 118.845 22.705 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 21.375 118.845 21.945 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 29.735 118.845 30.305 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 26.695 118.845 27.265 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 25.935 118.845 26.505 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 3.895 118.845 4.465 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 4.655 118.845 5.225 ;
  END
 END i18
 PIN i19
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 6.175 118.845 6.745 ;
  END
 END i19
 PIN i20
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 6.935 118.845 7.505 ;
  END
 END i20
 PIN i21
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 7.695 118.845 8.265 ;
  END
 END i21
 PIN i22
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 8.455 118.845 9.025 ;
  END
 END i22
 PIN i23
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 9.215 118.845 9.785 ;
  END
 END i23
 PIN i24
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 10.735 118.845 11.305 ;
  END
 END i24
 PIN i25
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 11.495 118.845 12.065 ;
  END
 END i25
 PIN i26
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 12.255 118.845 12.825 ;
  END
 END i26
 PIN i27
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 13.015 118.845 13.585 ;
  END
 END i27
 PIN i28
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 13.775 118.845 14.345 ;
  END
 END i28
 PIN i29
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 15.295 118.845 15.865 ;
  END
 END i29
 PIN i30
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 16.055 118.845 16.625 ;
  END
 END i30
 PIN i31
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 16.815 118.845 17.385 ;
  END
 END i31
 PIN i32
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 17.575 118.845 18.145 ;
  END
 END i32
 PIN i33
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 118.275 18.335 118.845 18.905 ;
  END
 END i33
 OBS
  LAYER metal1 ;
   RECT 0 0 121.98 61.56 ;
  LAYER via1 ;
   RECT 0 0 121.98 61.56 ;
  LAYER metal2 ;
   RECT 0 0 121.98 61.56 ;
  LAYER via2 ;
   RECT 0 0 121.98 61.56 ;
  LAYER metal3 ;
   RECT 0 0 121.98 61.56 ;
  LAYER via3 ;
   RECT 0 0 121.98 61.56 ;
  LAYER metal4 ;
   RECT 0 0 121.98 61.56 ;
 END
END block_321x324_65

MACRO block_779x1557_110
 CLASS BLOCK ;
 FOREIGN block_779x1557_110 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 296.02 BY 295.83 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 285.665 27.265 286.235 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 269.325 27.265 269.895 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 75.905 27.265 76.475 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 41.325 27.265 41.895 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 24.985 27.265 25.555 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 8.645 27.265 9.215 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 252.985 27.265 253.555 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 236.645 27.265 237.215 ;
  END
 END o7
 PIN o8
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 202.065 27.265 202.635 ;
  END
 END o8
 PIN o9
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 185.725 27.265 186.295 ;
  END
 END o9
 PIN o10
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 169.385 27.265 169.955 ;
  END
 END o10
 PIN o11
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 153.045 27.265 153.615 ;
  END
 END o11
 PIN o12
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 108.585 27.265 109.155 ;
  END
 END o12
 PIN o13
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 92.245 27.265 92.815 ;
  END
 END o13
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 142.025 4.085 142.595 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 124.925 4.085 125.495 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 136.705 4.085 137.275 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 132.335 4.085 132.905 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 129.485 4.085 130.055 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 4.275 141.645 4.845 142.215 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 4.275 142.405 4.845 142.975 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 142.785 4.085 143.355 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 133.095 4.085 133.665 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 119.985 4.085 120.555 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 4.275 125.305 4.845 125.875 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 128.535 4.085 129.105 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 125.685 4.085 126.255 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 123.595 4.085 124.165 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 121.125 4.085 121.695 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 4.275 119.605 4.845 120.175 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 13.015 143.165 13.585 143.735 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 13.015 129.865 13.585 130.435 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 287.375 27.265 287.945 ;
  END
 END i18
 PIN i19
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 271.035 27.265 271.605 ;
  END
 END i19
 PIN i20
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 74.195 27.265 74.765 ;
  END
 END i20
 PIN i21
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 39.615 27.265 40.185 ;
  END
 END i21
 PIN i22
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 23.275 27.265 23.845 ;
  END
 END i22
 PIN i23
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 6.935 27.265 7.505 ;
  END
 END i23
 PIN i24
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 254.695 27.265 255.265 ;
  END
 END i24
 PIN i25
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 238.355 27.265 238.925 ;
  END
 END i25
 PIN i26
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 203.775 27.265 204.345 ;
  END
 END i26
 PIN i27
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 187.435 27.265 188.005 ;
  END
 END i27
 PIN i28
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 171.095 27.265 171.665 ;
  END
 END i28
 PIN i29
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 154.755 27.265 155.325 ;
  END
 END i29
 PIN i30
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 106.875 27.265 107.445 ;
  END
 END i30
 PIN i31
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 90.535 27.265 91.105 ;
  END
 END i31
 PIN i32
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.455 252.415 28.025 252.985 ;
  END
 END i32
 PIN i33
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 248.425 27.265 248.995 ;
  END
 END i33
 PIN i34
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 244.245 27.265 244.815 ;
  END
 END i34
 PIN i35
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 260.585 27.265 261.155 ;
  END
 END i35
 PIN i36
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.455 185.155 28.025 185.725 ;
  END
 END i36
 PIN i37
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 181.165 27.265 181.735 ;
  END
 END i37
 PIN i38
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 176.985 27.265 177.555 ;
  END
 END i38
 PIN i39
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 172.995 27.265 173.565 ;
  END
 END i39
 PIN i40
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.455 92.815 28.025 93.385 ;
  END
 END i40
 PIN i41
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 96.805 27.265 97.375 ;
  END
 END i41
 PIN i42
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 100.985 27.265 101.555 ;
  END
 END i42
 PIN i43
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 104.975 27.265 105.545 ;
  END
 END i43
 PIN i44
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.455 25.555 28.025 26.125 ;
  END
 END i44
 PIN i45
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 29.545 27.265 30.115 ;
  END
 END i45
 PIN i46
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 33.725 27.265 34.295 ;
  END
 END i46
 PIN i47
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 17.385 27.265 17.955 ;
  END
 END i47
 PIN i48
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 256.595 27.265 257.165 ;
  END
 END i48
 PIN i49
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 189.335 27.265 189.905 ;
  END
 END i49
 PIN i50
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 88.635 27.265 89.205 ;
  END
 END i50
 PIN i51
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.695 21.375 27.265 21.945 ;
  END
 END i51
 PIN i52
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 18.335 143.165 18.905 143.735 ;
  END
 END i52
 PIN i53
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 18.335 129.865 18.905 130.435 ;
  END
 END i53
 PIN i54
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.455 286.805 28.025 287.375 ;
  END
 END i54
 PIN i55
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.455 270.465 28.025 271.035 ;
  END
 END i55
 PIN i56
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.455 74.765 28.025 75.335 ;
  END
 END i56
 PIN i57
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.455 40.185 28.025 40.755 ;
  END
 END i57
 PIN i58
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.455 23.845 28.025 24.415 ;
  END
 END i58
 PIN i59
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.455 7.505 28.025 8.075 ;
  END
 END i59
 PIN i60
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.455 254.125 28.025 254.695 ;
  END
 END i60
 PIN i61
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.455 237.785 28.025 238.355 ;
  END
 END i61
 PIN i62
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.455 203.205 28.025 203.775 ;
  END
 END i62
 PIN i63
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.455 186.865 28.025 187.435 ;
  END
 END i63
 PIN i64
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.455 170.525 28.025 171.095 ;
  END
 END i64
 PIN i65
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.455 154.185 28.025 154.755 ;
  END
 END i65
 PIN i66
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.455 107.445 28.025 108.015 ;
  END
 END i66
 PIN i67
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.455 91.105 28.025 91.675 ;
  END
 END i67
 PIN i68
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 135.565 4.085 136.135 ;
  END
 END i68
 PIN i69
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 4.275 135.185 4.845 135.755 ;
  END
 END i69
 PIN i70
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.215 286.235 28.785 286.805 ;
  END
 END i70
 PIN i71
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.215 269.895 28.785 270.465 ;
  END
 END i71
 PIN i72
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.215 75.335 28.785 75.905 ;
  END
 END i72
 PIN i73
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.215 40.755 28.785 41.325 ;
  END
 END i73
 PIN i74
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.215 24.415 28.785 24.985 ;
  END
 END i74
 PIN i75
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.215 8.075 28.785 8.645 ;
  END
 END i75
 PIN i76
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.215 253.555 28.785 254.125 ;
  END
 END i76
 PIN i77
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.215 237.215 28.785 237.785 ;
  END
 END i77
 PIN i78
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.215 202.635 28.785 203.205 ;
  END
 END i78
 PIN i79
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.215 186.295 28.785 186.865 ;
  END
 END i79
 PIN i80
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.215 169.955 28.785 170.525 ;
  END
 END i80
 PIN i81
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.215 153.615 28.785 154.185 ;
  END
 END i81
 PIN i82
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.215 108.015 28.785 108.585 ;
  END
 END i82
 PIN i83
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.215 91.675 28.785 92.245 ;
  END
 END i83
 PIN i84
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 4.275 143.165 4.845 143.735 ;
  END
 END i84
 PIN i85
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 5.415 143.165 5.985 143.735 ;
  END
 END i85
 PIN i86
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 7.315 143.165 7.885 143.735 ;
  END
 END i86
 PIN i87
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 8.835 143.165 9.405 143.735 ;
  END
 END i87
 PIN i88
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 143.165 10.925 143.735 ;
  END
 END i88
 PIN i89
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 12.255 143.165 12.825 143.735 ;
  END
 END i89
 PIN i90
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 4.275 129.865 4.845 130.435 ;
  END
 END i90
 PIN i91
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 5.415 129.865 5.985 130.435 ;
  END
 END i91
 PIN i92
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 7.315 129.865 7.885 130.435 ;
  END
 END i92
 PIN i93
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 8.835 129.865 9.405 130.435 ;
  END
 END i93
 PIN i94
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 129.865 10.925 130.435 ;
  END
 END i94
 PIN i95
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 12.255 129.865 12.825 130.435 ;
  END
 END i95
 OBS
  LAYER metal1 ;
   RECT 23.18 0.0 296.02 1.71 ;
   RECT 23.18 1.71 296.02 3.42 ;
   RECT 23.18 3.42 296.02 5.13 ;
   RECT 23.18 5.13 296.02 6.84 ;
   RECT 23.18 6.84 296.02 8.55 ;
   RECT 23.18 8.55 296.02 10.26 ;
   RECT 23.18 10.26 296.02 11.97 ;
   RECT 23.18 11.97 296.02 13.68 ;
   RECT 23.18 13.68 296.02 15.39 ;
   RECT 23.18 15.39 296.02 17.1 ;
   RECT 23.18 17.1 296.02 18.81 ;
   RECT 23.18 18.81 296.02 20.52 ;
   RECT 23.18 20.52 296.02 22.23 ;
   RECT 23.18 22.23 296.02 23.94 ;
   RECT 23.18 23.94 296.02 25.65 ;
   RECT 23.18 25.65 296.02 27.36 ;
   RECT 23.18 27.36 296.02 29.07 ;
   RECT 23.18 29.07 296.02 30.78 ;
   RECT 23.18 30.78 296.02 32.49 ;
   RECT 23.18 32.49 296.02 34.2 ;
   RECT 23.18 34.2 296.02 35.91 ;
   RECT 23.18 35.91 296.02 37.62 ;
   RECT 23.18 37.62 296.02 39.33 ;
   RECT 23.18 39.33 296.02 41.04 ;
   RECT 23.18 41.04 296.02 42.75 ;
   RECT 23.18 42.75 296.02 44.46 ;
   RECT 23.18 44.46 296.02 46.17 ;
   RECT 23.18 46.17 296.02 47.88 ;
   RECT 23.18 47.88 296.02 49.59 ;
   RECT 23.18 49.59 296.02 51.3 ;
   RECT 23.18 51.3 296.02 53.01 ;
   RECT 23.18 53.01 296.02 54.72 ;
   RECT 23.18 54.72 296.02 56.43 ;
   RECT 23.18 56.43 296.02 58.14 ;
   RECT 23.18 58.14 296.02 59.85 ;
   RECT 23.18 59.85 296.02 61.56 ;
   RECT 23.18 61.56 296.02 63.27 ;
   RECT 23.18 63.27 296.02 64.98 ;
   RECT 23.18 64.98 296.02 66.69 ;
   RECT 23.18 66.69 296.02 68.4 ;
   RECT 23.18 68.4 296.02 70.11 ;
   RECT 23.18 70.11 296.02 71.82 ;
   RECT 23.18 71.82 296.02 73.53 ;
   RECT 23.18 73.53 296.02 75.24 ;
   RECT 23.18 75.24 296.02 76.95 ;
   RECT 23.18 76.95 296.02 78.66 ;
   RECT 23.18 78.66 296.02 80.37 ;
   RECT 23.18 80.37 296.02 82.08 ;
   RECT 23.18 82.08 296.02 83.79 ;
   RECT 23.18 83.79 296.02 85.5 ;
   RECT 23.18 85.5 296.02 87.21 ;
   RECT 23.18 87.21 296.02 88.92 ;
   RECT 23.18 88.92 296.02 90.63 ;
   RECT 23.18 90.63 296.02 92.34 ;
   RECT 23.18 92.34 296.02 94.05 ;
   RECT 23.18 94.05 296.02 95.76 ;
   RECT 23.18 95.76 296.02 97.47 ;
   RECT 23.18 97.47 296.02 99.18 ;
   RECT 23.18 99.18 296.02 100.89 ;
   RECT 23.18 100.89 296.02 102.6 ;
   RECT 23.18 102.6 296.02 104.31 ;
   RECT 23.18 104.31 296.02 106.02 ;
   RECT 23.18 106.02 296.02 107.73 ;
   RECT 23.18 107.73 296.02 109.44 ;
   RECT 23.18 109.44 296.02 111.15 ;
   RECT 23.18 111.15 296.02 112.86 ;
   RECT 23.18 112.86 296.02 114.57 ;
   RECT 23.18 114.57 296.02 116.28 ;
   RECT 0.0 116.28 296.02 117.99 ;
   RECT 0.0 117.99 296.02 119.7 ;
   RECT 0.0 119.7 296.02 121.41 ;
   RECT 0.0 121.41 296.02 123.12 ;
   RECT 0.0 123.12 296.02 124.83 ;
   RECT 0.0 124.83 296.02 126.54 ;
   RECT 0.0 126.54 296.02 128.25 ;
   RECT 0.0 128.25 296.02 129.96 ;
   RECT 0.0 129.96 296.02 131.67 ;
   RECT 0.0 131.67 296.02 133.38 ;
   RECT 0.0 133.38 296.02 135.09 ;
   RECT 0.0 135.09 296.02 136.8 ;
   RECT 0.0 136.8 296.02 138.51 ;
   RECT 0.0 138.51 296.02 140.22 ;
   RECT 0.0 140.22 296.02 141.93 ;
   RECT 0.0 141.93 296.02 143.64 ;
   RECT 0.0 143.64 296.02 145.35 ;
   RECT 23.18 145.35 296.02 147.06 ;
   RECT 23.18 147.06 296.02 148.77 ;
   RECT 23.18 148.77 296.02 150.48 ;
   RECT 23.18 150.48 296.02 152.19 ;
   RECT 23.18 152.19 296.02 153.9 ;
   RECT 23.18 153.9 296.02 155.61 ;
   RECT 23.18 155.61 296.02 157.32 ;
   RECT 23.18 157.32 296.02 159.03 ;
   RECT 23.18 159.03 296.02 160.74 ;
   RECT 23.18 160.74 296.02 162.45 ;
   RECT 23.18 162.45 296.02 164.16 ;
   RECT 23.18 164.16 296.02 165.87 ;
   RECT 23.18 165.87 296.02 167.58 ;
   RECT 23.18 167.58 296.02 169.29 ;
   RECT 23.18 169.29 296.02 171.0 ;
   RECT 23.18 171.0 296.02 172.71 ;
   RECT 23.18 172.71 296.02 174.42 ;
   RECT 23.18 174.42 296.02 176.13 ;
   RECT 23.18 176.13 296.02 177.84 ;
   RECT 23.18 177.84 296.02 179.55 ;
   RECT 23.18 179.55 296.02 181.26 ;
   RECT 23.18 181.26 296.02 182.97 ;
   RECT 23.18 182.97 296.02 184.68 ;
   RECT 23.18 184.68 296.02 186.39 ;
   RECT 23.18 186.39 296.02 188.1 ;
   RECT 23.18 188.1 296.02 189.81 ;
   RECT 23.18 189.81 296.02 191.52 ;
   RECT 23.18 191.52 296.02 193.23 ;
   RECT 23.18 193.23 296.02 194.94 ;
   RECT 23.18 194.94 296.02 196.65 ;
   RECT 23.18 196.65 296.02 198.36 ;
   RECT 23.18 198.36 296.02 200.07 ;
   RECT 23.18 200.07 296.02 201.78 ;
   RECT 23.18 201.78 296.02 203.49 ;
   RECT 23.18 203.49 296.02 205.2 ;
   RECT 23.18 205.2 296.02 206.91 ;
   RECT 23.18 206.91 296.02 208.62 ;
   RECT 23.18 208.62 296.02 210.33 ;
   RECT 23.18 210.33 296.02 212.04 ;
   RECT 23.18 212.04 296.02 213.75 ;
   RECT 23.18 213.75 296.02 215.46 ;
   RECT 23.18 215.46 296.02 217.17 ;
   RECT 23.18 217.17 296.02 218.88 ;
   RECT 23.18 218.88 296.02 220.59 ;
   RECT 23.18 220.59 296.02 222.3 ;
   RECT 23.18 222.3 296.02 224.01 ;
   RECT 23.18 224.01 296.02 225.72 ;
   RECT 23.18 225.72 296.02 227.43 ;
   RECT 23.18 227.43 296.02 229.14 ;
   RECT 23.18 229.14 296.02 230.85 ;
   RECT 23.18 230.85 296.02 232.56 ;
   RECT 23.18 232.56 296.02 234.27 ;
   RECT 23.18 234.27 296.02 235.98 ;
   RECT 23.18 235.98 296.02 237.69 ;
   RECT 23.18 237.69 296.02 239.4 ;
   RECT 23.18 239.4 296.02 241.11 ;
   RECT 23.18 241.11 296.02 242.82 ;
   RECT 23.18 242.82 296.02 244.53 ;
   RECT 23.18 244.53 296.02 246.24 ;
   RECT 23.18 246.24 296.02 247.95 ;
   RECT 23.18 247.95 296.02 249.66 ;
   RECT 23.18 249.66 296.02 251.37 ;
   RECT 23.18 251.37 296.02 253.08 ;
   RECT 23.18 253.08 296.02 254.79 ;
   RECT 23.18 254.79 296.02 256.5 ;
   RECT 23.18 256.5 296.02 258.21 ;
   RECT 23.18 258.21 296.02 259.92 ;
   RECT 23.18 259.92 296.02 261.63 ;
   RECT 23.18 261.63 296.02 263.34 ;
   RECT 23.18 263.34 296.02 265.05 ;
   RECT 23.18 265.05 296.02 266.76 ;
   RECT 23.18 266.76 296.02 268.47 ;
   RECT 23.18 268.47 296.02 270.18 ;
   RECT 23.18 270.18 296.02 271.89 ;
   RECT 23.18 271.89 296.02 273.6 ;
   RECT 23.18 273.6 296.02 275.31 ;
   RECT 23.18 275.31 296.02 277.02 ;
   RECT 23.18 277.02 296.02 278.73 ;
   RECT 23.18 278.73 296.02 280.44 ;
   RECT 23.18 280.44 296.02 282.15 ;
   RECT 23.18 282.15 296.02 283.86 ;
   RECT 23.18 283.86 296.02 285.57 ;
   RECT 23.18 285.57 296.02 287.28 ;
   RECT 23.18 287.28 296.02 288.99 ;
   RECT 23.18 288.99 296.02 290.7 ;
   RECT 23.18 290.7 296.02 292.41 ;
   RECT 23.18 292.41 296.02 294.12 ;
   RECT 23.18 294.12 296.02 295.83 ;
  LAYER via1 ;
   RECT 23.18 0.0 296.02 1.71 ;
   RECT 23.18 1.71 296.02 3.42 ;
   RECT 23.18 3.42 296.02 5.13 ;
   RECT 23.18 5.13 296.02 6.84 ;
   RECT 23.18 6.84 296.02 8.55 ;
   RECT 23.18 8.55 296.02 10.26 ;
   RECT 23.18 10.26 296.02 11.97 ;
   RECT 23.18 11.97 296.02 13.68 ;
   RECT 23.18 13.68 296.02 15.39 ;
   RECT 23.18 15.39 296.02 17.1 ;
   RECT 23.18 17.1 296.02 18.81 ;
   RECT 23.18 18.81 296.02 20.52 ;
   RECT 23.18 20.52 296.02 22.23 ;
   RECT 23.18 22.23 296.02 23.94 ;
   RECT 23.18 23.94 296.02 25.65 ;
   RECT 23.18 25.65 296.02 27.36 ;
   RECT 23.18 27.36 296.02 29.07 ;
   RECT 23.18 29.07 296.02 30.78 ;
   RECT 23.18 30.78 296.02 32.49 ;
   RECT 23.18 32.49 296.02 34.2 ;
   RECT 23.18 34.2 296.02 35.91 ;
   RECT 23.18 35.91 296.02 37.62 ;
   RECT 23.18 37.62 296.02 39.33 ;
   RECT 23.18 39.33 296.02 41.04 ;
   RECT 23.18 41.04 296.02 42.75 ;
   RECT 23.18 42.75 296.02 44.46 ;
   RECT 23.18 44.46 296.02 46.17 ;
   RECT 23.18 46.17 296.02 47.88 ;
   RECT 23.18 47.88 296.02 49.59 ;
   RECT 23.18 49.59 296.02 51.3 ;
   RECT 23.18 51.3 296.02 53.01 ;
   RECT 23.18 53.01 296.02 54.72 ;
   RECT 23.18 54.72 296.02 56.43 ;
   RECT 23.18 56.43 296.02 58.14 ;
   RECT 23.18 58.14 296.02 59.85 ;
   RECT 23.18 59.85 296.02 61.56 ;
   RECT 23.18 61.56 296.02 63.27 ;
   RECT 23.18 63.27 296.02 64.98 ;
   RECT 23.18 64.98 296.02 66.69 ;
   RECT 23.18 66.69 296.02 68.4 ;
   RECT 23.18 68.4 296.02 70.11 ;
   RECT 23.18 70.11 296.02 71.82 ;
   RECT 23.18 71.82 296.02 73.53 ;
   RECT 23.18 73.53 296.02 75.24 ;
   RECT 23.18 75.24 296.02 76.95 ;
   RECT 23.18 76.95 296.02 78.66 ;
   RECT 23.18 78.66 296.02 80.37 ;
   RECT 23.18 80.37 296.02 82.08 ;
   RECT 23.18 82.08 296.02 83.79 ;
   RECT 23.18 83.79 296.02 85.5 ;
   RECT 23.18 85.5 296.02 87.21 ;
   RECT 23.18 87.21 296.02 88.92 ;
   RECT 23.18 88.92 296.02 90.63 ;
   RECT 23.18 90.63 296.02 92.34 ;
   RECT 23.18 92.34 296.02 94.05 ;
   RECT 23.18 94.05 296.02 95.76 ;
   RECT 23.18 95.76 296.02 97.47 ;
   RECT 23.18 97.47 296.02 99.18 ;
   RECT 23.18 99.18 296.02 100.89 ;
   RECT 23.18 100.89 296.02 102.6 ;
   RECT 23.18 102.6 296.02 104.31 ;
   RECT 23.18 104.31 296.02 106.02 ;
   RECT 23.18 106.02 296.02 107.73 ;
   RECT 23.18 107.73 296.02 109.44 ;
   RECT 23.18 109.44 296.02 111.15 ;
   RECT 23.18 111.15 296.02 112.86 ;
   RECT 23.18 112.86 296.02 114.57 ;
   RECT 23.18 114.57 296.02 116.28 ;
   RECT 0.0 116.28 296.02 117.99 ;
   RECT 0.0 117.99 296.02 119.7 ;
   RECT 0.0 119.7 296.02 121.41 ;
   RECT 0.0 121.41 296.02 123.12 ;
   RECT 0.0 123.12 296.02 124.83 ;
   RECT 0.0 124.83 296.02 126.54 ;
   RECT 0.0 126.54 296.02 128.25 ;
   RECT 0.0 128.25 296.02 129.96 ;
   RECT 0.0 129.96 296.02 131.67 ;
   RECT 0.0 131.67 296.02 133.38 ;
   RECT 0.0 133.38 296.02 135.09 ;
   RECT 0.0 135.09 296.02 136.8 ;
   RECT 0.0 136.8 296.02 138.51 ;
   RECT 0.0 138.51 296.02 140.22 ;
   RECT 0.0 140.22 296.02 141.93 ;
   RECT 0.0 141.93 296.02 143.64 ;
   RECT 0.0 143.64 296.02 145.35 ;
   RECT 23.18 145.35 296.02 147.06 ;
   RECT 23.18 147.06 296.02 148.77 ;
   RECT 23.18 148.77 296.02 150.48 ;
   RECT 23.18 150.48 296.02 152.19 ;
   RECT 23.18 152.19 296.02 153.9 ;
   RECT 23.18 153.9 296.02 155.61 ;
   RECT 23.18 155.61 296.02 157.32 ;
   RECT 23.18 157.32 296.02 159.03 ;
   RECT 23.18 159.03 296.02 160.74 ;
   RECT 23.18 160.74 296.02 162.45 ;
   RECT 23.18 162.45 296.02 164.16 ;
   RECT 23.18 164.16 296.02 165.87 ;
   RECT 23.18 165.87 296.02 167.58 ;
   RECT 23.18 167.58 296.02 169.29 ;
   RECT 23.18 169.29 296.02 171.0 ;
   RECT 23.18 171.0 296.02 172.71 ;
   RECT 23.18 172.71 296.02 174.42 ;
   RECT 23.18 174.42 296.02 176.13 ;
   RECT 23.18 176.13 296.02 177.84 ;
   RECT 23.18 177.84 296.02 179.55 ;
   RECT 23.18 179.55 296.02 181.26 ;
   RECT 23.18 181.26 296.02 182.97 ;
   RECT 23.18 182.97 296.02 184.68 ;
   RECT 23.18 184.68 296.02 186.39 ;
   RECT 23.18 186.39 296.02 188.1 ;
   RECT 23.18 188.1 296.02 189.81 ;
   RECT 23.18 189.81 296.02 191.52 ;
   RECT 23.18 191.52 296.02 193.23 ;
   RECT 23.18 193.23 296.02 194.94 ;
   RECT 23.18 194.94 296.02 196.65 ;
   RECT 23.18 196.65 296.02 198.36 ;
   RECT 23.18 198.36 296.02 200.07 ;
   RECT 23.18 200.07 296.02 201.78 ;
   RECT 23.18 201.78 296.02 203.49 ;
   RECT 23.18 203.49 296.02 205.2 ;
   RECT 23.18 205.2 296.02 206.91 ;
   RECT 23.18 206.91 296.02 208.62 ;
   RECT 23.18 208.62 296.02 210.33 ;
   RECT 23.18 210.33 296.02 212.04 ;
   RECT 23.18 212.04 296.02 213.75 ;
   RECT 23.18 213.75 296.02 215.46 ;
   RECT 23.18 215.46 296.02 217.17 ;
   RECT 23.18 217.17 296.02 218.88 ;
   RECT 23.18 218.88 296.02 220.59 ;
   RECT 23.18 220.59 296.02 222.3 ;
   RECT 23.18 222.3 296.02 224.01 ;
   RECT 23.18 224.01 296.02 225.72 ;
   RECT 23.18 225.72 296.02 227.43 ;
   RECT 23.18 227.43 296.02 229.14 ;
   RECT 23.18 229.14 296.02 230.85 ;
   RECT 23.18 230.85 296.02 232.56 ;
   RECT 23.18 232.56 296.02 234.27 ;
   RECT 23.18 234.27 296.02 235.98 ;
   RECT 23.18 235.98 296.02 237.69 ;
   RECT 23.18 237.69 296.02 239.4 ;
   RECT 23.18 239.4 296.02 241.11 ;
   RECT 23.18 241.11 296.02 242.82 ;
   RECT 23.18 242.82 296.02 244.53 ;
   RECT 23.18 244.53 296.02 246.24 ;
   RECT 23.18 246.24 296.02 247.95 ;
   RECT 23.18 247.95 296.02 249.66 ;
   RECT 23.18 249.66 296.02 251.37 ;
   RECT 23.18 251.37 296.02 253.08 ;
   RECT 23.18 253.08 296.02 254.79 ;
   RECT 23.18 254.79 296.02 256.5 ;
   RECT 23.18 256.5 296.02 258.21 ;
   RECT 23.18 258.21 296.02 259.92 ;
   RECT 23.18 259.92 296.02 261.63 ;
   RECT 23.18 261.63 296.02 263.34 ;
   RECT 23.18 263.34 296.02 265.05 ;
   RECT 23.18 265.05 296.02 266.76 ;
   RECT 23.18 266.76 296.02 268.47 ;
   RECT 23.18 268.47 296.02 270.18 ;
   RECT 23.18 270.18 296.02 271.89 ;
   RECT 23.18 271.89 296.02 273.6 ;
   RECT 23.18 273.6 296.02 275.31 ;
   RECT 23.18 275.31 296.02 277.02 ;
   RECT 23.18 277.02 296.02 278.73 ;
   RECT 23.18 278.73 296.02 280.44 ;
   RECT 23.18 280.44 296.02 282.15 ;
   RECT 23.18 282.15 296.02 283.86 ;
   RECT 23.18 283.86 296.02 285.57 ;
   RECT 23.18 285.57 296.02 287.28 ;
   RECT 23.18 287.28 296.02 288.99 ;
   RECT 23.18 288.99 296.02 290.7 ;
   RECT 23.18 290.7 296.02 292.41 ;
   RECT 23.18 292.41 296.02 294.12 ;
   RECT 23.18 294.12 296.02 295.83 ;
  LAYER metal2 ;
   RECT 23.18 0.0 296.02 1.71 ;
   RECT 23.18 1.71 296.02 3.42 ;
   RECT 23.18 3.42 296.02 5.13 ;
   RECT 23.18 5.13 296.02 6.84 ;
   RECT 23.18 6.84 296.02 8.55 ;
   RECT 23.18 8.55 296.02 10.26 ;
   RECT 23.18 10.26 296.02 11.97 ;
   RECT 23.18 11.97 296.02 13.68 ;
   RECT 23.18 13.68 296.02 15.39 ;
   RECT 23.18 15.39 296.02 17.1 ;
   RECT 23.18 17.1 296.02 18.81 ;
   RECT 23.18 18.81 296.02 20.52 ;
   RECT 23.18 20.52 296.02 22.23 ;
   RECT 23.18 22.23 296.02 23.94 ;
   RECT 23.18 23.94 296.02 25.65 ;
   RECT 23.18 25.65 296.02 27.36 ;
   RECT 23.18 27.36 296.02 29.07 ;
   RECT 23.18 29.07 296.02 30.78 ;
   RECT 23.18 30.78 296.02 32.49 ;
   RECT 23.18 32.49 296.02 34.2 ;
   RECT 23.18 34.2 296.02 35.91 ;
   RECT 23.18 35.91 296.02 37.62 ;
   RECT 23.18 37.62 296.02 39.33 ;
   RECT 23.18 39.33 296.02 41.04 ;
   RECT 23.18 41.04 296.02 42.75 ;
   RECT 23.18 42.75 296.02 44.46 ;
   RECT 23.18 44.46 296.02 46.17 ;
   RECT 23.18 46.17 296.02 47.88 ;
   RECT 23.18 47.88 296.02 49.59 ;
   RECT 23.18 49.59 296.02 51.3 ;
   RECT 23.18 51.3 296.02 53.01 ;
   RECT 23.18 53.01 296.02 54.72 ;
   RECT 23.18 54.72 296.02 56.43 ;
   RECT 23.18 56.43 296.02 58.14 ;
   RECT 23.18 58.14 296.02 59.85 ;
   RECT 23.18 59.85 296.02 61.56 ;
   RECT 23.18 61.56 296.02 63.27 ;
   RECT 23.18 63.27 296.02 64.98 ;
   RECT 23.18 64.98 296.02 66.69 ;
   RECT 23.18 66.69 296.02 68.4 ;
   RECT 23.18 68.4 296.02 70.11 ;
   RECT 23.18 70.11 296.02 71.82 ;
   RECT 23.18 71.82 296.02 73.53 ;
   RECT 23.18 73.53 296.02 75.24 ;
   RECT 23.18 75.24 296.02 76.95 ;
   RECT 23.18 76.95 296.02 78.66 ;
   RECT 23.18 78.66 296.02 80.37 ;
   RECT 23.18 80.37 296.02 82.08 ;
   RECT 23.18 82.08 296.02 83.79 ;
   RECT 23.18 83.79 296.02 85.5 ;
   RECT 23.18 85.5 296.02 87.21 ;
   RECT 23.18 87.21 296.02 88.92 ;
   RECT 23.18 88.92 296.02 90.63 ;
   RECT 23.18 90.63 296.02 92.34 ;
   RECT 23.18 92.34 296.02 94.05 ;
   RECT 23.18 94.05 296.02 95.76 ;
   RECT 23.18 95.76 296.02 97.47 ;
   RECT 23.18 97.47 296.02 99.18 ;
   RECT 23.18 99.18 296.02 100.89 ;
   RECT 23.18 100.89 296.02 102.6 ;
   RECT 23.18 102.6 296.02 104.31 ;
   RECT 23.18 104.31 296.02 106.02 ;
   RECT 23.18 106.02 296.02 107.73 ;
   RECT 23.18 107.73 296.02 109.44 ;
   RECT 23.18 109.44 296.02 111.15 ;
   RECT 23.18 111.15 296.02 112.86 ;
   RECT 23.18 112.86 296.02 114.57 ;
   RECT 23.18 114.57 296.02 116.28 ;
   RECT 0.0 116.28 296.02 117.99 ;
   RECT 0.0 117.99 296.02 119.7 ;
   RECT 0.0 119.7 296.02 121.41 ;
   RECT 0.0 121.41 296.02 123.12 ;
   RECT 0.0 123.12 296.02 124.83 ;
   RECT 0.0 124.83 296.02 126.54 ;
   RECT 0.0 126.54 296.02 128.25 ;
   RECT 0.0 128.25 296.02 129.96 ;
   RECT 0.0 129.96 296.02 131.67 ;
   RECT 0.0 131.67 296.02 133.38 ;
   RECT 0.0 133.38 296.02 135.09 ;
   RECT 0.0 135.09 296.02 136.8 ;
   RECT 0.0 136.8 296.02 138.51 ;
   RECT 0.0 138.51 296.02 140.22 ;
   RECT 0.0 140.22 296.02 141.93 ;
   RECT 0.0 141.93 296.02 143.64 ;
   RECT 0.0 143.64 296.02 145.35 ;
   RECT 23.18 145.35 296.02 147.06 ;
   RECT 23.18 147.06 296.02 148.77 ;
   RECT 23.18 148.77 296.02 150.48 ;
   RECT 23.18 150.48 296.02 152.19 ;
   RECT 23.18 152.19 296.02 153.9 ;
   RECT 23.18 153.9 296.02 155.61 ;
   RECT 23.18 155.61 296.02 157.32 ;
   RECT 23.18 157.32 296.02 159.03 ;
   RECT 23.18 159.03 296.02 160.74 ;
   RECT 23.18 160.74 296.02 162.45 ;
   RECT 23.18 162.45 296.02 164.16 ;
   RECT 23.18 164.16 296.02 165.87 ;
   RECT 23.18 165.87 296.02 167.58 ;
   RECT 23.18 167.58 296.02 169.29 ;
   RECT 23.18 169.29 296.02 171.0 ;
   RECT 23.18 171.0 296.02 172.71 ;
   RECT 23.18 172.71 296.02 174.42 ;
   RECT 23.18 174.42 296.02 176.13 ;
   RECT 23.18 176.13 296.02 177.84 ;
   RECT 23.18 177.84 296.02 179.55 ;
   RECT 23.18 179.55 296.02 181.26 ;
   RECT 23.18 181.26 296.02 182.97 ;
   RECT 23.18 182.97 296.02 184.68 ;
   RECT 23.18 184.68 296.02 186.39 ;
   RECT 23.18 186.39 296.02 188.1 ;
   RECT 23.18 188.1 296.02 189.81 ;
   RECT 23.18 189.81 296.02 191.52 ;
   RECT 23.18 191.52 296.02 193.23 ;
   RECT 23.18 193.23 296.02 194.94 ;
   RECT 23.18 194.94 296.02 196.65 ;
   RECT 23.18 196.65 296.02 198.36 ;
   RECT 23.18 198.36 296.02 200.07 ;
   RECT 23.18 200.07 296.02 201.78 ;
   RECT 23.18 201.78 296.02 203.49 ;
   RECT 23.18 203.49 296.02 205.2 ;
   RECT 23.18 205.2 296.02 206.91 ;
   RECT 23.18 206.91 296.02 208.62 ;
   RECT 23.18 208.62 296.02 210.33 ;
   RECT 23.18 210.33 296.02 212.04 ;
   RECT 23.18 212.04 296.02 213.75 ;
   RECT 23.18 213.75 296.02 215.46 ;
   RECT 23.18 215.46 296.02 217.17 ;
   RECT 23.18 217.17 296.02 218.88 ;
   RECT 23.18 218.88 296.02 220.59 ;
   RECT 23.18 220.59 296.02 222.3 ;
   RECT 23.18 222.3 296.02 224.01 ;
   RECT 23.18 224.01 296.02 225.72 ;
   RECT 23.18 225.72 296.02 227.43 ;
   RECT 23.18 227.43 296.02 229.14 ;
   RECT 23.18 229.14 296.02 230.85 ;
   RECT 23.18 230.85 296.02 232.56 ;
   RECT 23.18 232.56 296.02 234.27 ;
   RECT 23.18 234.27 296.02 235.98 ;
   RECT 23.18 235.98 296.02 237.69 ;
   RECT 23.18 237.69 296.02 239.4 ;
   RECT 23.18 239.4 296.02 241.11 ;
   RECT 23.18 241.11 296.02 242.82 ;
   RECT 23.18 242.82 296.02 244.53 ;
   RECT 23.18 244.53 296.02 246.24 ;
   RECT 23.18 246.24 296.02 247.95 ;
   RECT 23.18 247.95 296.02 249.66 ;
   RECT 23.18 249.66 296.02 251.37 ;
   RECT 23.18 251.37 296.02 253.08 ;
   RECT 23.18 253.08 296.02 254.79 ;
   RECT 23.18 254.79 296.02 256.5 ;
   RECT 23.18 256.5 296.02 258.21 ;
   RECT 23.18 258.21 296.02 259.92 ;
   RECT 23.18 259.92 296.02 261.63 ;
   RECT 23.18 261.63 296.02 263.34 ;
   RECT 23.18 263.34 296.02 265.05 ;
   RECT 23.18 265.05 296.02 266.76 ;
   RECT 23.18 266.76 296.02 268.47 ;
   RECT 23.18 268.47 296.02 270.18 ;
   RECT 23.18 270.18 296.02 271.89 ;
   RECT 23.18 271.89 296.02 273.6 ;
   RECT 23.18 273.6 296.02 275.31 ;
   RECT 23.18 275.31 296.02 277.02 ;
   RECT 23.18 277.02 296.02 278.73 ;
   RECT 23.18 278.73 296.02 280.44 ;
   RECT 23.18 280.44 296.02 282.15 ;
   RECT 23.18 282.15 296.02 283.86 ;
   RECT 23.18 283.86 296.02 285.57 ;
   RECT 23.18 285.57 296.02 287.28 ;
   RECT 23.18 287.28 296.02 288.99 ;
   RECT 23.18 288.99 296.02 290.7 ;
   RECT 23.18 290.7 296.02 292.41 ;
   RECT 23.18 292.41 296.02 294.12 ;
   RECT 23.18 294.12 296.02 295.83 ;
  LAYER via2 ;
   RECT 23.18 0.0 296.02 1.71 ;
   RECT 23.18 1.71 296.02 3.42 ;
   RECT 23.18 3.42 296.02 5.13 ;
   RECT 23.18 5.13 296.02 6.84 ;
   RECT 23.18 6.84 296.02 8.55 ;
   RECT 23.18 8.55 296.02 10.26 ;
   RECT 23.18 10.26 296.02 11.97 ;
   RECT 23.18 11.97 296.02 13.68 ;
   RECT 23.18 13.68 296.02 15.39 ;
   RECT 23.18 15.39 296.02 17.1 ;
   RECT 23.18 17.1 296.02 18.81 ;
   RECT 23.18 18.81 296.02 20.52 ;
   RECT 23.18 20.52 296.02 22.23 ;
   RECT 23.18 22.23 296.02 23.94 ;
   RECT 23.18 23.94 296.02 25.65 ;
   RECT 23.18 25.65 296.02 27.36 ;
   RECT 23.18 27.36 296.02 29.07 ;
   RECT 23.18 29.07 296.02 30.78 ;
   RECT 23.18 30.78 296.02 32.49 ;
   RECT 23.18 32.49 296.02 34.2 ;
   RECT 23.18 34.2 296.02 35.91 ;
   RECT 23.18 35.91 296.02 37.62 ;
   RECT 23.18 37.62 296.02 39.33 ;
   RECT 23.18 39.33 296.02 41.04 ;
   RECT 23.18 41.04 296.02 42.75 ;
   RECT 23.18 42.75 296.02 44.46 ;
   RECT 23.18 44.46 296.02 46.17 ;
   RECT 23.18 46.17 296.02 47.88 ;
   RECT 23.18 47.88 296.02 49.59 ;
   RECT 23.18 49.59 296.02 51.3 ;
   RECT 23.18 51.3 296.02 53.01 ;
   RECT 23.18 53.01 296.02 54.72 ;
   RECT 23.18 54.72 296.02 56.43 ;
   RECT 23.18 56.43 296.02 58.14 ;
   RECT 23.18 58.14 296.02 59.85 ;
   RECT 23.18 59.85 296.02 61.56 ;
   RECT 23.18 61.56 296.02 63.27 ;
   RECT 23.18 63.27 296.02 64.98 ;
   RECT 23.18 64.98 296.02 66.69 ;
   RECT 23.18 66.69 296.02 68.4 ;
   RECT 23.18 68.4 296.02 70.11 ;
   RECT 23.18 70.11 296.02 71.82 ;
   RECT 23.18 71.82 296.02 73.53 ;
   RECT 23.18 73.53 296.02 75.24 ;
   RECT 23.18 75.24 296.02 76.95 ;
   RECT 23.18 76.95 296.02 78.66 ;
   RECT 23.18 78.66 296.02 80.37 ;
   RECT 23.18 80.37 296.02 82.08 ;
   RECT 23.18 82.08 296.02 83.79 ;
   RECT 23.18 83.79 296.02 85.5 ;
   RECT 23.18 85.5 296.02 87.21 ;
   RECT 23.18 87.21 296.02 88.92 ;
   RECT 23.18 88.92 296.02 90.63 ;
   RECT 23.18 90.63 296.02 92.34 ;
   RECT 23.18 92.34 296.02 94.05 ;
   RECT 23.18 94.05 296.02 95.76 ;
   RECT 23.18 95.76 296.02 97.47 ;
   RECT 23.18 97.47 296.02 99.18 ;
   RECT 23.18 99.18 296.02 100.89 ;
   RECT 23.18 100.89 296.02 102.6 ;
   RECT 23.18 102.6 296.02 104.31 ;
   RECT 23.18 104.31 296.02 106.02 ;
   RECT 23.18 106.02 296.02 107.73 ;
   RECT 23.18 107.73 296.02 109.44 ;
   RECT 23.18 109.44 296.02 111.15 ;
   RECT 23.18 111.15 296.02 112.86 ;
   RECT 23.18 112.86 296.02 114.57 ;
   RECT 23.18 114.57 296.02 116.28 ;
   RECT 0.0 116.28 296.02 117.99 ;
   RECT 0.0 117.99 296.02 119.7 ;
   RECT 0.0 119.7 296.02 121.41 ;
   RECT 0.0 121.41 296.02 123.12 ;
   RECT 0.0 123.12 296.02 124.83 ;
   RECT 0.0 124.83 296.02 126.54 ;
   RECT 0.0 126.54 296.02 128.25 ;
   RECT 0.0 128.25 296.02 129.96 ;
   RECT 0.0 129.96 296.02 131.67 ;
   RECT 0.0 131.67 296.02 133.38 ;
   RECT 0.0 133.38 296.02 135.09 ;
   RECT 0.0 135.09 296.02 136.8 ;
   RECT 0.0 136.8 296.02 138.51 ;
   RECT 0.0 138.51 296.02 140.22 ;
   RECT 0.0 140.22 296.02 141.93 ;
   RECT 0.0 141.93 296.02 143.64 ;
   RECT 0.0 143.64 296.02 145.35 ;
   RECT 23.18 145.35 296.02 147.06 ;
   RECT 23.18 147.06 296.02 148.77 ;
   RECT 23.18 148.77 296.02 150.48 ;
   RECT 23.18 150.48 296.02 152.19 ;
   RECT 23.18 152.19 296.02 153.9 ;
   RECT 23.18 153.9 296.02 155.61 ;
   RECT 23.18 155.61 296.02 157.32 ;
   RECT 23.18 157.32 296.02 159.03 ;
   RECT 23.18 159.03 296.02 160.74 ;
   RECT 23.18 160.74 296.02 162.45 ;
   RECT 23.18 162.45 296.02 164.16 ;
   RECT 23.18 164.16 296.02 165.87 ;
   RECT 23.18 165.87 296.02 167.58 ;
   RECT 23.18 167.58 296.02 169.29 ;
   RECT 23.18 169.29 296.02 171.0 ;
   RECT 23.18 171.0 296.02 172.71 ;
   RECT 23.18 172.71 296.02 174.42 ;
   RECT 23.18 174.42 296.02 176.13 ;
   RECT 23.18 176.13 296.02 177.84 ;
   RECT 23.18 177.84 296.02 179.55 ;
   RECT 23.18 179.55 296.02 181.26 ;
   RECT 23.18 181.26 296.02 182.97 ;
   RECT 23.18 182.97 296.02 184.68 ;
   RECT 23.18 184.68 296.02 186.39 ;
   RECT 23.18 186.39 296.02 188.1 ;
   RECT 23.18 188.1 296.02 189.81 ;
   RECT 23.18 189.81 296.02 191.52 ;
   RECT 23.18 191.52 296.02 193.23 ;
   RECT 23.18 193.23 296.02 194.94 ;
   RECT 23.18 194.94 296.02 196.65 ;
   RECT 23.18 196.65 296.02 198.36 ;
   RECT 23.18 198.36 296.02 200.07 ;
   RECT 23.18 200.07 296.02 201.78 ;
   RECT 23.18 201.78 296.02 203.49 ;
   RECT 23.18 203.49 296.02 205.2 ;
   RECT 23.18 205.2 296.02 206.91 ;
   RECT 23.18 206.91 296.02 208.62 ;
   RECT 23.18 208.62 296.02 210.33 ;
   RECT 23.18 210.33 296.02 212.04 ;
   RECT 23.18 212.04 296.02 213.75 ;
   RECT 23.18 213.75 296.02 215.46 ;
   RECT 23.18 215.46 296.02 217.17 ;
   RECT 23.18 217.17 296.02 218.88 ;
   RECT 23.18 218.88 296.02 220.59 ;
   RECT 23.18 220.59 296.02 222.3 ;
   RECT 23.18 222.3 296.02 224.01 ;
   RECT 23.18 224.01 296.02 225.72 ;
   RECT 23.18 225.72 296.02 227.43 ;
   RECT 23.18 227.43 296.02 229.14 ;
   RECT 23.18 229.14 296.02 230.85 ;
   RECT 23.18 230.85 296.02 232.56 ;
   RECT 23.18 232.56 296.02 234.27 ;
   RECT 23.18 234.27 296.02 235.98 ;
   RECT 23.18 235.98 296.02 237.69 ;
   RECT 23.18 237.69 296.02 239.4 ;
   RECT 23.18 239.4 296.02 241.11 ;
   RECT 23.18 241.11 296.02 242.82 ;
   RECT 23.18 242.82 296.02 244.53 ;
   RECT 23.18 244.53 296.02 246.24 ;
   RECT 23.18 246.24 296.02 247.95 ;
   RECT 23.18 247.95 296.02 249.66 ;
   RECT 23.18 249.66 296.02 251.37 ;
   RECT 23.18 251.37 296.02 253.08 ;
   RECT 23.18 253.08 296.02 254.79 ;
   RECT 23.18 254.79 296.02 256.5 ;
   RECT 23.18 256.5 296.02 258.21 ;
   RECT 23.18 258.21 296.02 259.92 ;
   RECT 23.18 259.92 296.02 261.63 ;
   RECT 23.18 261.63 296.02 263.34 ;
   RECT 23.18 263.34 296.02 265.05 ;
   RECT 23.18 265.05 296.02 266.76 ;
   RECT 23.18 266.76 296.02 268.47 ;
   RECT 23.18 268.47 296.02 270.18 ;
   RECT 23.18 270.18 296.02 271.89 ;
   RECT 23.18 271.89 296.02 273.6 ;
   RECT 23.18 273.6 296.02 275.31 ;
   RECT 23.18 275.31 296.02 277.02 ;
   RECT 23.18 277.02 296.02 278.73 ;
   RECT 23.18 278.73 296.02 280.44 ;
   RECT 23.18 280.44 296.02 282.15 ;
   RECT 23.18 282.15 296.02 283.86 ;
   RECT 23.18 283.86 296.02 285.57 ;
   RECT 23.18 285.57 296.02 287.28 ;
   RECT 23.18 287.28 296.02 288.99 ;
   RECT 23.18 288.99 296.02 290.7 ;
   RECT 23.18 290.7 296.02 292.41 ;
   RECT 23.18 292.41 296.02 294.12 ;
   RECT 23.18 294.12 296.02 295.83 ;
  LAYER metal3 ;
   RECT 23.18 0.0 296.02 1.71 ;
   RECT 23.18 1.71 296.02 3.42 ;
   RECT 23.18 3.42 296.02 5.13 ;
   RECT 23.18 5.13 296.02 6.84 ;
   RECT 23.18 6.84 296.02 8.55 ;
   RECT 23.18 8.55 296.02 10.26 ;
   RECT 23.18 10.26 296.02 11.97 ;
   RECT 23.18 11.97 296.02 13.68 ;
   RECT 23.18 13.68 296.02 15.39 ;
   RECT 23.18 15.39 296.02 17.1 ;
   RECT 23.18 17.1 296.02 18.81 ;
   RECT 23.18 18.81 296.02 20.52 ;
   RECT 23.18 20.52 296.02 22.23 ;
   RECT 23.18 22.23 296.02 23.94 ;
   RECT 23.18 23.94 296.02 25.65 ;
   RECT 23.18 25.65 296.02 27.36 ;
   RECT 23.18 27.36 296.02 29.07 ;
   RECT 23.18 29.07 296.02 30.78 ;
   RECT 23.18 30.78 296.02 32.49 ;
   RECT 23.18 32.49 296.02 34.2 ;
   RECT 23.18 34.2 296.02 35.91 ;
   RECT 23.18 35.91 296.02 37.62 ;
   RECT 23.18 37.62 296.02 39.33 ;
   RECT 23.18 39.33 296.02 41.04 ;
   RECT 23.18 41.04 296.02 42.75 ;
   RECT 23.18 42.75 296.02 44.46 ;
   RECT 23.18 44.46 296.02 46.17 ;
   RECT 23.18 46.17 296.02 47.88 ;
   RECT 23.18 47.88 296.02 49.59 ;
   RECT 23.18 49.59 296.02 51.3 ;
   RECT 23.18 51.3 296.02 53.01 ;
   RECT 23.18 53.01 296.02 54.72 ;
   RECT 23.18 54.72 296.02 56.43 ;
   RECT 23.18 56.43 296.02 58.14 ;
   RECT 23.18 58.14 296.02 59.85 ;
   RECT 23.18 59.85 296.02 61.56 ;
   RECT 23.18 61.56 296.02 63.27 ;
   RECT 23.18 63.27 296.02 64.98 ;
   RECT 23.18 64.98 296.02 66.69 ;
   RECT 23.18 66.69 296.02 68.4 ;
   RECT 23.18 68.4 296.02 70.11 ;
   RECT 23.18 70.11 296.02 71.82 ;
   RECT 23.18 71.82 296.02 73.53 ;
   RECT 23.18 73.53 296.02 75.24 ;
   RECT 23.18 75.24 296.02 76.95 ;
   RECT 23.18 76.95 296.02 78.66 ;
   RECT 23.18 78.66 296.02 80.37 ;
   RECT 23.18 80.37 296.02 82.08 ;
   RECT 23.18 82.08 296.02 83.79 ;
   RECT 23.18 83.79 296.02 85.5 ;
   RECT 23.18 85.5 296.02 87.21 ;
   RECT 23.18 87.21 296.02 88.92 ;
   RECT 23.18 88.92 296.02 90.63 ;
   RECT 23.18 90.63 296.02 92.34 ;
   RECT 23.18 92.34 296.02 94.05 ;
   RECT 23.18 94.05 296.02 95.76 ;
   RECT 23.18 95.76 296.02 97.47 ;
   RECT 23.18 97.47 296.02 99.18 ;
   RECT 23.18 99.18 296.02 100.89 ;
   RECT 23.18 100.89 296.02 102.6 ;
   RECT 23.18 102.6 296.02 104.31 ;
   RECT 23.18 104.31 296.02 106.02 ;
   RECT 23.18 106.02 296.02 107.73 ;
   RECT 23.18 107.73 296.02 109.44 ;
   RECT 23.18 109.44 296.02 111.15 ;
   RECT 23.18 111.15 296.02 112.86 ;
   RECT 23.18 112.86 296.02 114.57 ;
   RECT 23.18 114.57 296.02 116.28 ;
   RECT 0.0 116.28 296.02 117.99 ;
   RECT 0.0 117.99 296.02 119.7 ;
   RECT 0.0 119.7 296.02 121.41 ;
   RECT 0.0 121.41 296.02 123.12 ;
   RECT 0.0 123.12 296.02 124.83 ;
   RECT 0.0 124.83 296.02 126.54 ;
   RECT 0.0 126.54 296.02 128.25 ;
   RECT 0.0 128.25 296.02 129.96 ;
   RECT 0.0 129.96 296.02 131.67 ;
   RECT 0.0 131.67 296.02 133.38 ;
   RECT 0.0 133.38 296.02 135.09 ;
   RECT 0.0 135.09 296.02 136.8 ;
   RECT 0.0 136.8 296.02 138.51 ;
   RECT 0.0 138.51 296.02 140.22 ;
   RECT 0.0 140.22 296.02 141.93 ;
   RECT 0.0 141.93 296.02 143.64 ;
   RECT 0.0 143.64 296.02 145.35 ;
   RECT 23.18 145.35 296.02 147.06 ;
   RECT 23.18 147.06 296.02 148.77 ;
   RECT 23.18 148.77 296.02 150.48 ;
   RECT 23.18 150.48 296.02 152.19 ;
   RECT 23.18 152.19 296.02 153.9 ;
   RECT 23.18 153.9 296.02 155.61 ;
   RECT 23.18 155.61 296.02 157.32 ;
   RECT 23.18 157.32 296.02 159.03 ;
   RECT 23.18 159.03 296.02 160.74 ;
   RECT 23.18 160.74 296.02 162.45 ;
   RECT 23.18 162.45 296.02 164.16 ;
   RECT 23.18 164.16 296.02 165.87 ;
   RECT 23.18 165.87 296.02 167.58 ;
   RECT 23.18 167.58 296.02 169.29 ;
   RECT 23.18 169.29 296.02 171.0 ;
   RECT 23.18 171.0 296.02 172.71 ;
   RECT 23.18 172.71 296.02 174.42 ;
   RECT 23.18 174.42 296.02 176.13 ;
   RECT 23.18 176.13 296.02 177.84 ;
   RECT 23.18 177.84 296.02 179.55 ;
   RECT 23.18 179.55 296.02 181.26 ;
   RECT 23.18 181.26 296.02 182.97 ;
   RECT 23.18 182.97 296.02 184.68 ;
   RECT 23.18 184.68 296.02 186.39 ;
   RECT 23.18 186.39 296.02 188.1 ;
   RECT 23.18 188.1 296.02 189.81 ;
   RECT 23.18 189.81 296.02 191.52 ;
   RECT 23.18 191.52 296.02 193.23 ;
   RECT 23.18 193.23 296.02 194.94 ;
   RECT 23.18 194.94 296.02 196.65 ;
   RECT 23.18 196.65 296.02 198.36 ;
   RECT 23.18 198.36 296.02 200.07 ;
   RECT 23.18 200.07 296.02 201.78 ;
   RECT 23.18 201.78 296.02 203.49 ;
   RECT 23.18 203.49 296.02 205.2 ;
   RECT 23.18 205.2 296.02 206.91 ;
   RECT 23.18 206.91 296.02 208.62 ;
   RECT 23.18 208.62 296.02 210.33 ;
   RECT 23.18 210.33 296.02 212.04 ;
   RECT 23.18 212.04 296.02 213.75 ;
   RECT 23.18 213.75 296.02 215.46 ;
   RECT 23.18 215.46 296.02 217.17 ;
   RECT 23.18 217.17 296.02 218.88 ;
   RECT 23.18 218.88 296.02 220.59 ;
   RECT 23.18 220.59 296.02 222.3 ;
   RECT 23.18 222.3 296.02 224.01 ;
   RECT 23.18 224.01 296.02 225.72 ;
   RECT 23.18 225.72 296.02 227.43 ;
   RECT 23.18 227.43 296.02 229.14 ;
   RECT 23.18 229.14 296.02 230.85 ;
   RECT 23.18 230.85 296.02 232.56 ;
   RECT 23.18 232.56 296.02 234.27 ;
   RECT 23.18 234.27 296.02 235.98 ;
   RECT 23.18 235.98 296.02 237.69 ;
   RECT 23.18 237.69 296.02 239.4 ;
   RECT 23.18 239.4 296.02 241.11 ;
   RECT 23.18 241.11 296.02 242.82 ;
   RECT 23.18 242.82 296.02 244.53 ;
   RECT 23.18 244.53 296.02 246.24 ;
   RECT 23.18 246.24 296.02 247.95 ;
   RECT 23.18 247.95 296.02 249.66 ;
   RECT 23.18 249.66 296.02 251.37 ;
   RECT 23.18 251.37 296.02 253.08 ;
   RECT 23.18 253.08 296.02 254.79 ;
   RECT 23.18 254.79 296.02 256.5 ;
   RECT 23.18 256.5 296.02 258.21 ;
   RECT 23.18 258.21 296.02 259.92 ;
   RECT 23.18 259.92 296.02 261.63 ;
   RECT 23.18 261.63 296.02 263.34 ;
   RECT 23.18 263.34 296.02 265.05 ;
   RECT 23.18 265.05 296.02 266.76 ;
   RECT 23.18 266.76 296.02 268.47 ;
   RECT 23.18 268.47 296.02 270.18 ;
   RECT 23.18 270.18 296.02 271.89 ;
   RECT 23.18 271.89 296.02 273.6 ;
   RECT 23.18 273.6 296.02 275.31 ;
   RECT 23.18 275.31 296.02 277.02 ;
   RECT 23.18 277.02 296.02 278.73 ;
   RECT 23.18 278.73 296.02 280.44 ;
   RECT 23.18 280.44 296.02 282.15 ;
   RECT 23.18 282.15 296.02 283.86 ;
   RECT 23.18 283.86 296.02 285.57 ;
   RECT 23.18 285.57 296.02 287.28 ;
   RECT 23.18 287.28 296.02 288.99 ;
   RECT 23.18 288.99 296.02 290.7 ;
   RECT 23.18 290.7 296.02 292.41 ;
   RECT 23.18 292.41 296.02 294.12 ;
   RECT 23.18 294.12 296.02 295.83 ;
  LAYER via3 ;
   RECT 23.18 0.0 296.02 1.71 ;
   RECT 23.18 1.71 296.02 3.42 ;
   RECT 23.18 3.42 296.02 5.13 ;
   RECT 23.18 5.13 296.02 6.84 ;
   RECT 23.18 6.84 296.02 8.55 ;
   RECT 23.18 8.55 296.02 10.26 ;
   RECT 23.18 10.26 296.02 11.97 ;
   RECT 23.18 11.97 296.02 13.68 ;
   RECT 23.18 13.68 296.02 15.39 ;
   RECT 23.18 15.39 296.02 17.1 ;
   RECT 23.18 17.1 296.02 18.81 ;
   RECT 23.18 18.81 296.02 20.52 ;
   RECT 23.18 20.52 296.02 22.23 ;
   RECT 23.18 22.23 296.02 23.94 ;
   RECT 23.18 23.94 296.02 25.65 ;
   RECT 23.18 25.65 296.02 27.36 ;
   RECT 23.18 27.36 296.02 29.07 ;
   RECT 23.18 29.07 296.02 30.78 ;
   RECT 23.18 30.78 296.02 32.49 ;
   RECT 23.18 32.49 296.02 34.2 ;
   RECT 23.18 34.2 296.02 35.91 ;
   RECT 23.18 35.91 296.02 37.62 ;
   RECT 23.18 37.62 296.02 39.33 ;
   RECT 23.18 39.33 296.02 41.04 ;
   RECT 23.18 41.04 296.02 42.75 ;
   RECT 23.18 42.75 296.02 44.46 ;
   RECT 23.18 44.46 296.02 46.17 ;
   RECT 23.18 46.17 296.02 47.88 ;
   RECT 23.18 47.88 296.02 49.59 ;
   RECT 23.18 49.59 296.02 51.3 ;
   RECT 23.18 51.3 296.02 53.01 ;
   RECT 23.18 53.01 296.02 54.72 ;
   RECT 23.18 54.72 296.02 56.43 ;
   RECT 23.18 56.43 296.02 58.14 ;
   RECT 23.18 58.14 296.02 59.85 ;
   RECT 23.18 59.85 296.02 61.56 ;
   RECT 23.18 61.56 296.02 63.27 ;
   RECT 23.18 63.27 296.02 64.98 ;
   RECT 23.18 64.98 296.02 66.69 ;
   RECT 23.18 66.69 296.02 68.4 ;
   RECT 23.18 68.4 296.02 70.11 ;
   RECT 23.18 70.11 296.02 71.82 ;
   RECT 23.18 71.82 296.02 73.53 ;
   RECT 23.18 73.53 296.02 75.24 ;
   RECT 23.18 75.24 296.02 76.95 ;
   RECT 23.18 76.95 296.02 78.66 ;
   RECT 23.18 78.66 296.02 80.37 ;
   RECT 23.18 80.37 296.02 82.08 ;
   RECT 23.18 82.08 296.02 83.79 ;
   RECT 23.18 83.79 296.02 85.5 ;
   RECT 23.18 85.5 296.02 87.21 ;
   RECT 23.18 87.21 296.02 88.92 ;
   RECT 23.18 88.92 296.02 90.63 ;
   RECT 23.18 90.63 296.02 92.34 ;
   RECT 23.18 92.34 296.02 94.05 ;
   RECT 23.18 94.05 296.02 95.76 ;
   RECT 23.18 95.76 296.02 97.47 ;
   RECT 23.18 97.47 296.02 99.18 ;
   RECT 23.18 99.18 296.02 100.89 ;
   RECT 23.18 100.89 296.02 102.6 ;
   RECT 23.18 102.6 296.02 104.31 ;
   RECT 23.18 104.31 296.02 106.02 ;
   RECT 23.18 106.02 296.02 107.73 ;
   RECT 23.18 107.73 296.02 109.44 ;
   RECT 23.18 109.44 296.02 111.15 ;
   RECT 23.18 111.15 296.02 112.86 ;
   RECT 23.18 112.86 296.02 114.57 ;
   RECT 23.18 114.57 296.02 116.28 ;
   RECT 0.0 116.28 296.02 117.99 ;
   RECT 0.0 117.99 296.02 119.7 ;
   RECT 0.0 119.7 296.02 121.41 ;
   RECT 0.0 121.41 296.02 123.12 ;
   RECT 0.0 123.12 296.02 124.83 ;
   RECT 0.0 124.83 296.02 126.54 ;
   RECT 0.0 126.54 296.02 128.25 ;
   RECT 0.0 128.25 296.02 129.96 ;
   RECT 0.0 129.96 296.02 131.67 ;
   RECT 0.0 131.67 296.02 133.38 ;
   RECT 0.0 133.38 296.02 135.09 ;
   RECT 0.0 135.09 296.02 136.8 ;
   RECT 0.0 136.8 296.02 138.51 ;
   RECT 0.0 138.51 296.02 140.22 ;
   RECT 0.0 140.22 296.02 141.93 ;
   RECT 0.0 141.93 296.02 143.64 ;
   RECT 0.0 143.64 296.02 145.35 ;
   RECT 23.18 145.35 296.02 147.06 ;
   RECT 23.18 147.06 296.02 148.77 ;
   RECT 23.18 148.77 296.02 150.48 ;
   RECT 23.18 150.48 296.02 152.19 ;
   RECT 23.18 152.19 296.02 153.9 ;
   RECT 23.18 153.9 296.02 155.61 ;
   RECT 23.18 155.61 296.02 157.32 ;
   RECT 23.18 157.32 296.02 159.03 ;
   RECT 23.18 159.03 296.02 160.74 ;
   RECT 23.18 160.74 296.02 162.45 ;
   RECT 23.18 162.45 296.02 164.16 ;
   RECT 23.18 164.16 296.02 165.87 ;
   RECT 23.18 165.87 296.02 167.58 ;
   RECT 23.18 167.58 296.02 169.29 ;
   RECT 23.18 169.29 296.02 171.0 ;
   RECT 23.18 171.0 296.02 172.71 ;
   RECT 23.18 172.71 296.02 174.42 ;
   RECT 23.18 174.42 296.02 176.13 ;
   RECT 23.18 176.13 296.02 177.84 ;
   RECT 23.18 177.84 296.02 179.55 ;
   RECT 23.18 179.55 296.02 181.26 ;
   RECT 23.18 181.26 296.02 182.97 ;
   RECT 23.18 182.97 296.02 184.68 ;
   RECT 23.18 184.68 296.02 186.39 ;
   RECT 23.18 186.39 296.02 188.1 ;
   RECT 23.18 188.1 296.02 189.81 ;
   RECT 23.18 189.81 296.02 191.52 ;
   RECT 23.18 191.52 296.02 193.23 ;
   RECT 23.18 193.23 296.02 194.94 ;
   RECT 23.18 194.94 296.02 196.65 ;
   RECT 23.18 196.65 296.02 198.36 ;
   RECT 23.18 198.36 296.02 200.07 ;
   RECT 23.18 200.07 296.02 201.78 ;
   RECT 23.18 201.78 296.02 203.49 ;
   RECT 23.18 203.49 296.02 205.2 ;
   RECT 23.18 205.2 296.02 206.91 ;
   RECT 23.18 206.91 296.02 208.62 ;
   RECT 23.18 208.62 296.02 210.33 ;
   RECT 23.18 210.33 296.02 212.04 ;
   RECT 23.18 212.04 296.02 213.75 ;
   RECT 23.18 213.75 296.02 215.46 ;
   RECT 23.18 215.46 296.02 217.17 ;
   RECT 23.18 217.17 296.02 218.88 ;
   RECT 23.18 218.88 296.02 220.59 ;
   RECT 23.18 220.59 296.02 222.3 ;
   RECT 23.18 222.3 296.02 224.01 ;
   RECT 23.18 224.01 296.02 225.72 ;
   RECT 23.18 225.72 296.02 227.43 ;
   RECT 23.18 227.43 296.02 229.14 ;
   RECT 23.18 229.14 296.02 230.85 ;
   RECT 23.18 230.85 296.02 232.56 ;
   RECT 23.18 232.56 296.02 234.27 ;
   RECT 23.18 234.27 296.02 235.98 ;
   RECT 23.18 235.98 296.02 237.69 ;
   RECT 23.18 237.69 296.02 239.4 ;
   RECT 23.18 239.4 296.02 241.11 ;
   RECT 23.18 241.11 296.02 242.82 ;
   RECT 23.18 242.82 296.02 244.53 ;
   RECT 23.18 244.53 296.02 246.24 ;
   RECT 23.18 246.24 296.02 247.95 ;
   RECT 23.18 247.95 296.02 249.66 ;
   RECT 23.18 249.66 296.02 251.37 ;
   RECT 23.18 251.37 296.02 253.08 ;
   RECT 23.18 253.08 296.02 254.79 ;
   RECT 23.18 254.79 296.02 256.5 ;
   RECT 23.18 256.5 296.02 258.21 ;
   RECT 23.18 258.21 296.02 259.92 ;
   RECT 23.18 259.92 296.02 261.63 ;
   RECT 23.18 261.63 296.02 263.34 ;
   RECT 23.18 263.34 296.02 265.05 ;
   RECT 23.18 265.05 296.02 266.76 ;
   RECT 23.18 266.76 296.02 268.47 ;
   RECT 23.18 268.47 296.02 270.18 ;
   RECT 23.18 270.18 296.02 271.89 ;
   RECT 23.18 271.89 296.02 273.6 ;
   RECT 23.18 273.6 296.02 275.31 ;
   RECT 23.18 275.31 296.02 277.02 ;
   RECT 23.18 277.02 296.02 278.73 ;
   RECT 23.18 278.73 296.02 280.44 ;
   RECT 23.18 280.44 296.02 282.15 ;
   RECT 23.18 282.15 296.02 283.86 ;
   RECT 23.18 283.86 296.02 285.57 ;
   RECT 23.18 285.57 296.02 287.28 ;
   RECT 23.18 287.28 296.02 288.99 ;
   RECT 23.18 288.99 296.02 290.7 ;
   RECT 23.18 290.7 296.02 292.41 ;
   RECT 23.18 292.41 296.02 294.12 ;
   RECT 23.18 294.12 296.02 295.83 ;
  LAYER metal4 ;
   RECT 23.18 0.0 296.02 1.71 ;
   RECT 23.18 1.71 296.02 3.42 ;
   RECT 23.18 3.42 296.02 5.13 ;
   RECT 23.18 5.13 296.02 6.84 ;
   RECT 23.18 6.84 296.02 8.55 ;
   RECT 23.18 8.55 296.02 10.26 ;
   RECT 23.18 10.26 296.02 11.97 ;
   RECT 23.18 11.97 296.02 13.68 ;
   RECT 23.18 13.68 296.02 15.39 ;
   RECT 23.18 15.39 296.02 17.1 ;
   RECT 23.18 17.1 296.02 18.81 ;
   RECT 23.18 18.81 296.02 20.52 ;
   RECT 23.18 20.52 296.02 22.23 ;
   RECT 23.18 22.23 296.02 23.94 ;
   RECT 23.18 23.94 296.02 25.65 ;
   RECT 23.18 25.65 296.02 27.36 ;
   RECT 23.18 27.36 296.02 29.07 ;
   RECT 23.18 29.07 296.02 30.78 ;
   RECT 23.18 30.78 296.02 32.49 ;
   RECT 23.18 32.49 296.02 34.2 ;
   RECT 23.18 34.2 296.02 35.91 ;
   RECT 23.18 35.91 296.02 37.62 ;
   RECT 23.18 37.62 296.02 39.33 ;
   RECT 23.18 39.33 296.02 41.04 ;
   RECT 23.18 41.04 296.02 42.75 ;
   RECT 23.18 42.75 296.02 44.46 ;
   RECT 23.18 44.46 296.02 46.17 ;
   RECT 23.18 46.17 296.02 47.88 ;
   RECT 23.18 47.88 296.02 49.59 ;
   RECT 23.18 49.59 296.02 51.3 ;
   RECT 23.18 51.3 296.02 53.01 ;
   RECT 23.18 53.01 296.02 54.72 ;
   RECT 23.18 54.72 296.02 56.43 ;
   RECT 23.18 56.43 296.02 58.14 ;
   RECT 23.18 58.14 296.02 59.85 ;
   RECT 23.18 59.85 296.02 61.56 ;
   RECT 23.18 61.56 296.02 63.27 ;
   RECT 23.18 63.27 296.02 64.98 ;
   RECT 23.18 64.98 296.02 66.69 ;
   RECT 23.18 66.69 296.02 68.4 ;
   RECT 23.18 68.4 296.02 70.11 ;
   RECT 23.18 70.11 296.02 71.82 ;
   RECT 23.18 71.82 296.02 73.53 ;
   RECT 23.18 73.53 296.02 75.24 ;
   RECT 23.18 75.24 296.02 76.95 ;
   RECT 23.18 76.95 296.02 78.66 ;
   RECT 23.18 78.66 296.02 80.37 ;
   RECT 23.18 80.37 296.02 82.08 ;
   RECT 23.18 82.08 296.02 83.79 ;
   RECT 23.18 83.79 296.02 85.5 ;
   RECT 23.18 85.5 296.02 87.21 ;
   RECT 23.18 87.21 296.02 88.92 ;
   RECT 23.18 88.92 296.02 90.63 ;
   RECT 23.18 90.63 296.02 92.34 ;
   RECT 23.18 92.34 296.02 94.05 ;
   RECT 23.18 94.05 296.02 95.76 ;
   RECT 23.18 95.76 296.02 97.47 ;
   RECT 23.18 97.47 296.02 99.18 ;
   RECT 23.18 99.18 296.02 100.89 ;
   RECT 23.18 100.89 296.02 102.6 ;
   RECT 23.18 102.6 296.02 104.31 ;
   RECT 23.18 104.31 296.02 106.02 ;
   RECT 23.18 106.02 296.02 107.73 ;
   RECT 23.18 107.73 296.02 109.44 ;
   RECT 23.18 109.44 296.02 111.15 ;
   RECT 23.18 111.15 296.02 112.86 ;
   RECT 23.18 112.86 296.02 114.57 ;
   RECT 23.18 114.57 296.02 116.28 ;
   RECT 0.0 116.28 296.02 117.99 ;
   RECT 0.0 117.99 296.02 119.7 ;
   RECT 0.0 119.7 296.02 121.41 ;
   RECT 0.0 121.41 296.02 123.12 ;
   RECT 0.0 123.12 296.02 124.83 ;
   RECT 0.0 124.83 296.02 126.54 ;
   RECT 0.0 126.54 296.02 128.25 ;
   RECT 0.0 128.25 296.02 129.96 ;
   RECT 0.0 129.96 296.02 131.67 ;
   RECT 0.0 131.67 296.02 133.38 ;
   RECT 0.0 133.38 296.02 135.09 ;
   RECT 0.0 135.09 296.02 136.8 ;
   RECT 0.0 136.8 296.02 138.51 ;
   RECT 0.0 138.51 296.02 140.22 ;
   RECT 0.0 140.22 296.02 141.93 ;
   RECT 0.0 141.93 296.02 143.64 ;
   RECT 0.0 143.64 296.02 145.35 ;
   RECT 23.18 145.35 296.02 147.06 ;
   RECT 23.18 147.06 296.02 148.77 ;
   RECT 23.18 148.77 296.02 150.48 ;
   RECT 23.18 150.48 296.02 152.19 ;
   RECT 23.18 152.19 296.02 153.9 ;
   RECT 23.18 153.9 296.02 155.61 ;
   RECT 23.18 155.61 296.02 157.32 ;
   RECT 23.18 157.32 296.02 159.03 ;
   RECT 23.18 159.03 296.02 160.74 ;
   RECT 23.18 160.74 296.02 162.45 ;
   RECT 23.18 162.45 296.02 164.16 ;
   RECT 23.18 164.16 296.02 165.87 ;
   RECT 23.18 165.87 296.02 167.58 ;
   RECT 23.18 167.58 296.02 169.29 ;
   RECT 23.18 169.29 296.02 171.0 ;
   RECT 23.18 171.0 296.02 172.71 ;
   RECT 23.18 172.71 296.02 174.42 ;
   RECT 23.18 174.42 296.02 176.13 ;
   RECT 23.18 176.13 296.02 177.84 ;
   RECT 23.18 177.84 296.02 179.55 ;
   RECT 23.18 179.55 296.02 181.26 ;
   RECT 23.18 181.26 296.02 182.97 ;
   RECT 23.18 182.97 296.02 184.68 ;
   RECT 23.18 184.68 296.02 186.39 ;
   RECT 23.18 186.39 296.02 188.1 ;
   RECT 23.18 188.1 296.02 189.81 ;
   RECT 23.18 189.81 296.02 191.52 ;
   RECT 23.18 191.52 296.02 193.23 ;
   RECT 23.18 193.23 296.02 194.94 ;
   RECT 23.18 194.94 296.02 196.65 ;
   RECT 23.18 196.65 296.02 198.36 ;
   RECT 23.18 198.36 296.02 200.07 ;
   RECT 23.18 200.07 296.02 201.78 ;
   RECT 23.18 201.78 296.02 203.49 ;
   RECT 23.18 203.49 296.02 205.2 ;
   RECT 23.18 205.2 296.02 206.91 ;
   RECT 23.18 206.91 296.02 208.62 ;
   RECT 23.18 208.62 296.02 210.33 ;
   RECT 23.18 210.33 296.02 212.04 ;
   RECT 23.18 212.04 296.02 213.75 ;
   RECT 23.18 213.75 296.02 215.46 ;
   RECT 23.18 215.46 296.02 217.17 ;
   RECT 23.18 217.17 296.02 218.88 ;
   RECT 23.18 218.88 296.02 220.59 ;
   RECT 23.18 220.59 296.02 222.3 ;
   RECT 23.18 222.3 296.02 224.01 ;
   RECT 23.18 224.01 296.02 225.72 ;
   RECT 23.18 225.72 296.02 227.43 ;
   RECT 23.18 227.43 296.02 229.14 ;
   RECT 23.18 229.14 296.02 230.85 ;
   RECT 23.18 230.85 296.02 232.56 ;
   RECT 23.18 232.56 296.02 234.27 ;
   RECT 23.18 234.27 296.02 235.98 ;
   RECT 23.18 235.98 296.02 237.69 ;
   RECT 23.18 237.69 296.02 239.4 ;
   RECT 23.18 239.4 296.02 241.11 ;
   RECT 23.18 241.11 296.02 242.82 ;
   RECT 23.18 242.82 296.02 244.53 ;
   RECT 23.18 244.53 296.02 246.24 ;
   RECT 23.18 246.24 296.02 247.95 ;
   RECT 23.18 247.95 296.02 249.66 ;
   RECT 23.18 249.66 296.02 251.37 ;
   RECT 23.18 251.37 296.02 253.08 ;
   RECT 23.18 253.08 296.02 254.79 ;
   RECT 23.18 254.79 296.02 256.5 ;
   RECT 23.18 256.5 296.02 258.21 ;
   RECT 23.18 258.21 296.02 259.92 ;
   RECT 23.18 259.92 296.02 261.63 ;
   RECT 23.18 261.63 296.02 263.34 ;
   RECT 23.18 263.34 296.02 265.05 ;
   RECT 23.18 265.05 296.02 266.76 ;
   RECT 23.18 266.76 296.02 268.47 ;
   RECT 23.18 268.47 296.02 270.18 ;
   RECT 23.18 270.18 296.02 271.89 ;
   RECT 23.18 271.89 296.02 273.6 ;
   RECT 23.18 273.6 296.02 275.31 ;
   RECT 23.18 275.31 296.02 277.02 ;
   RECT 23.18 277.02 296.02 278.73 ;
   RECT 23.18 278.73 296.02 280.44 ;
   RECT 23.18 280.44 296.02 282.15 ;
   RECT 23.18 282.15 296.02 283.86 ;
   RECT 23.18 283.86 296.02 285.57 ;
   RECT 23.18 285.57 296.02 287.28 ;
   RECT 23.18 287.28 296.02 288.99 ;
   RECT 23.18 288.99 296.02 290.7 ;
   RECT 23.18 290.7 296.02 292.41 ;
   RECT 23.18 292.41 296.02 294.12 ;
   RECT 23.18 294.12 296.02 295.83 ;
 END
END block_779x1557_110

MACRO block_315x558_44
 CLASS BLOCK ;
 FOREIGN block_315x558_44 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 119.7 BY 106.02 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 102.885 9.785 103.455 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 19.665 9.785 20.235 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 13.965 9.785 14.535 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 8.265 9.785 8.835 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 2.375 9.785 2.945 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 97.185 9.785 97.755 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 91.485 9.785 92.055 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 85.785 9.785 86.355 ;
  END
 END o7
 PIN o8
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 79.895 9.785 80.465 ;
  END
 END o8
 PIN o9
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 74.195 9.785 74.765 ;
  END
 END o9
 PIN o10
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 68.495 9.785 69.065 ;
  END
 END o10
 PIN o11
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 36.955 9.785 37.525 ;
  END
 END o11
 PIN o12
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 31.255 9.785 31.825 ;
  END
 END o12
 PIN o13
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 25.365 9.785 25.935 ;
  END
 END o13
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 54.055 118.465 54.625 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 46.075 118.465 46.645 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 47.405 118.465 47.975 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 44.745 118.465 45.315 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.135 47.975 117.705 48.545 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 111.815 44.935 112.385 45.505 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 45.505 9.785 46.075 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 61.465 118.465 62.035 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 51.585 118.465 52.155 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 52.725 118.465 53.295 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 52.535 9.785 53.105 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 8.455 59.375 9.025 59.945 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 56.335 9.785 56.905 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.135 54.625 117.705 55.195 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 56.335 118.465 56.905 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.135 56.905 117.705 57.475 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 102.505 118.465 103.075 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 20.045 118.465 20.615 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 14.345 118.465 14.915 ;
  END
 END i18
 PIN i19
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 8.645 118.465 9.215 ;
  END
 END i19
 PIN i20
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 2.945 118.465 3.515 ;
  END
 END i20
 PIN i21
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 96.805 118.465 97.375 ;
  END
 END i21
 PIN i22
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 91.105 118.465 91.675 ;
  END
 END i22
 PIN i23
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 85.215 118.465 85.785 ;
  END
 END i23
 PIN i24
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 79.515 118.465 80.085 ;
  END
 END i24
 PIN i25
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 73.815 118.465 74.385 ;
  END
 END i25
 PIN i26
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 68.115 118.465 68.685 ;
  END
 END i26
 PIN i27
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 37.335 118.465 37.905 ;
  END
 END i27
 PIN i28
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 31.635 118.465 32.205 ;
  END
 END i28
 PIN i29
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 25.935 118.465 26.505 ;
  END
 END i29
 OBS
  LAYER metal1 ;
   RECT 0 0 119.7 106.02 ;
  LAYER via1 ;
   RECT 0 0 119.7 106.02 ;
  LAYER metal2 ;
   RECT 0 0 119.7 106.02 ;
  LAYER via2 ;
   RECT 0 0 119.7 106.02 ;
  LAYER metal3 ;
   RECT 0 0 119.7 106.02 ;
  LAYER via3 ;
   RECT 0 0 119.7 106.02 ;
  LAYER metal4 ;
   RECT 0 0 119.7 106.02 ;
 END
END block_315x558_44

MACRO block_414x3978_702
 CLASS BLOCK ;
 FOREIGN block_414x3978_702 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 157.32 BY 755.82 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 749.075 26.885 749.645 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 744.895 26.885 745.465 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 708.225 26.885 708.795 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 256.595 26.885 257.165 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 252.415 26.885 252.985 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 248.425 26.885 248.995 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 244.245 26.885 244.815 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 240.255 26.885 240.825 ;
  END
 END o7
 PIN o8
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 236.075 26.885 236.645 ;
  END
 END o8
 PIN o9
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 232.085 26.885 232.655 ;
  END
 END o9
 PIN o10
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 227.905 26.885 228.475 ;
  END
 END o10
 PIN o11
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 223.915 26.885 224.485 ;
  END
 END o11
 PIN o12
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 219.735 26.885 220.305 ;
  END
 END o12
 PIN o13
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 704.045 26.885 704.615 ;
  END
 END o13
 PIN o14
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 215.745 26.885 216.315 ;
  END
 END o14
 PIN o15
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 211.565 26.885 212.135 ;
  END
 END o15
 PIN o16
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 207.575 26.885 208.145 ;
  END
 END o16
 PIN o17
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 203.395 26.885 203.965 ;
  END
 END o17
 PIN o18
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 199.405 26.885 199.975 ;
  END
 END o18
 PIN o19
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 195.225 26.885 195.795 ;
  END
 END o19
 PIN o20
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 191.235 26.885 191.805 ;
  END
 END o20
 PIN o21
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 187.055 26.885 187.625 ;
  END
 END o21
 PIN o22
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 183.065 26.885 183.635 ;
  END
 END o22
 PIN o23
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 173.755 26.885 174.325 ;
  END
 END o23
 PIN o24
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 700.055 26.885 700.625 ;
  END
 END o24
 PIN o25
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 169.765 26.885 170.335 ;
  END
 END o25
 PIN o26
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 165.585 26.885 166.155 ;
  END
 END o26
 PIN o27
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 161.595 26.885 162.165 ;
  END
 END o27
 PIN o28
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 157.415 26.885 157.985 ;
  END
 END o28
 PIN o29
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 153.425 26.885 153.995 ;
  END
 END o29
 PIN o30
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 149.245 26.885 149.815 ;
  END
 END o30
 PIN o31
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 145.255 26.885 145.825 ;
  END
 END o31
 PIN o32
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 141.075 26.885 141.645 ;
  END
 END o32
 PIN o33
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 137.085 26.885 137.655 ;
  END
 END o33
 PIN o34
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 132.905 26.885 133.475 ;
  END
 END o34
 PIN o35
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 695.875 26.885 696.445 ;
  END
 END o35
 PIN o36
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 128.915 26.885 129.485 ;
  END
 END o36
 PIN o37
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 124.735 26.885 125.305 ;
  END
 END o37
 PIN o38
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 120.745 26.885 121.315 ;
  END
 END o38
 PIN o39
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 116.565 26.885 117.135 ;
  END
 END o39
 PIN o40
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 112.575 26.885 113.145 ;
  END
 END o40
 PIN o41
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 108.395 26.885 108.965 ;
  END
 END o41
 PIN o42
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 104.405 26.885 104.975 ;
  END
 END o42
 PIN o43
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 100.225 26.885 100.795 ;
  END
 END o43
 PIN o44
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 77.995 26.885 78.565 ;
  END
 END o44
 PIN o45
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 73.815 26.885 74.385 ;
  END
 END o45
 PIN o46
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 691.885 26.885 692.455 ;
  END
 END o46
 PIN o47
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 69.825 26.885 70.395 ;
  END
 END o47
 PIN o48
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 65.645 26.885 66.215 ;
  END
 END o48
 PIN o49
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 61.655 26.885 62.225 ;
  END
 END o49
 PIN o50
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 57.475 26.885 58.045 ;
  END
 END o50
 PIN o51
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 53.485 26.885 54.055 ;
  END
 END o51
 PIN o52
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 49.305 26.885 49.875 ;
  END
 END o52
 PIN o53
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 45.315 26.885 45.885 ;
  END
 END o53
 PIN o54
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 41.135 26.885 41.705 ;
  END
 END o54
 PIN o55
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 37.145 26.885 37.715 ;
  END
 END o55
 PIN o56
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 32.965 26.885 33.535 ;
  END
 END o56
 PIN o57
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 687.705 26.885 688.275 ;
  END
 END o57
 PIN o58
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 28.975 26.885 29.545 ;
  END
 END o58
 PIN o59
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 24.795 26.885 25.365 ;
  END
 END o59
 PIN o60
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 20.805 26.885 21.375 ;
  END
 END o60
 PIN o61
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 16.625 26.885 17.195 ;
  END
 END o61
 PIN o62
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 12.635 26.885 13.205 ;
  END
 END o62
 PIN o63
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 8.455 26.885 9.025 ;
  END
 END o63
 PIN o64
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 4.465 26.885 5.035 ;
  END
 END o64
 PIN o65
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 683.715 26.885 684.285 ;
  END
 END o65
 PIN o66
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 679.535 26.885 680.105 ;
  END
 END o66
 PIN o67
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 675.545 26.885 676.115 ;
  END
 END o67
 PIN o68
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 671.365 26.885 671.935 ;
  END
 END o68
 PIN o69
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 740.905 26.885 741.475 ;
  END
 END o69
 PIN o70
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 649.135 26.885 649.705 ;
  END
 END o70
 PIN o71
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 644.955 26.885 645.525 ;
  END
 END o71
 PIN o72
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 640.965 26.885 641.535 ;
  END
 END o72
 PIN o73
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 636.785 26.885 637.355 ;
  END
 END o73
 PIN o74
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 632.795 26.885 633.365 ;
  END
 END o74
 PIN o75
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 628.615 26.885 629.185 ;
  END
 END o75
 PIN o76
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 624.625 26.885 625.195 ;
  END
 END o76
 PIN o77
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 620.445 26.885 621.015 ;
  END
 END o77
 PIN o78
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 616.455 26.885 617.025 ;
  END
 END o78
 PIN o79
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 612.275 26.885 612.845 ;
  END
 END o79
 PIN o80
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 736.725 26.885 737.295 ;
  END
 END o80
 PIN o81
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 608.285 26.885 608.855 ;
  END
 END o81
 PIN o82
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 604.105 26.885 604.675 ;
  END
 END o82
 PIN o83
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 600.115 26.885 600.685 ;
  END
 END o83
 PIN o84
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 595.935 26.885 596.505 ;
  END
 END o84
 PIN o85
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 591.945 26.885 592.515 ;
  END
 END o85
 PIN o86
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 587.765 26.885 588.335 ;
  END
 END o86
 PIN o87
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 583.775 26.885 584.345 ;
  END
 END o87
 PIN o88
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 579.595 26.885 580.165 ;
  END
 END o88
 PIN o89
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 575.605 26.885 576.175 ;
  END
 END o89
 PIN o90
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 571.425 26.885 571.995 ;
  END
 END o90
 PIN o91
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 732.735 26.885 733.305 ;
  END
 END o91
 PIN o92
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 562.305 26.885 562.875 ;
  END
 END o92
 PIN o93
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 558.125 26.885 558.695 ;
  END
 END o93
 PIN o94
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 554.135 26.885 554.705 ;
  END
 END o94
 PIN o95
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 549.955 26.885 550.525 ;
  END
 END o95
 PIN o96
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 545.965 26.885 546.535 ;
  END
 END o96
 PIN o97
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 541.785 26.885 542.355 ;
  END
 END o97
 PIN o98
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 537.795 26.885 538.365 ;
  END
 END o98
 PIN o99
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 533.615 26.885 534.185 ;
  END
 END o99
 PIN o100
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 529.625 26.885 530.195 ;
  END
 END o100
 PIN o101
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 525.445 26.885 526.015 ;
  END
 END o101
 PIN o102
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 728.555 26.885 729.125 ;
  END
 END o102
 PIN o103
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 521.455 26.885 522.025 ;
  END
 END o103
 PIN o104
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 517.275 26.885 517.845 ;
  END
 END o104
 PIN o105
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 513.285 26.885 513.855 ;
  END
 END o105
 PIN o106
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 509.105 26.885 509.675 ;
  END
 END o106
 PIN o107
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 505.115 26.885 505.685 ;
  END
 END o107
 PIN o108
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 500.935 26.885 501.505 ;
  END
 END o108
 PIN o109
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 496.945 26.885 497.515 ;
  END
 END o109
 PIN o110
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 492.765 26.885 493.335 ;
  END
 END o110
 PIN o111
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 488.775 26.885 489.345 ;
  END
 END o111
 PIN o112
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 484.595 26.885 485.165 ;
  END
 END o112
 PIN o113
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 724.565 26.885 725.135 ;
  END
 END o113
 PIN o114
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 462.365 26.885 462.935 ;
  END
 END o114
 PIN o115
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 458.185 26.885 458.755 ;
  END
 END o115
 PIN o116
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 454.195 26.885 454.765 ;
  END
 END o116
 PIN o117
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 450.015 26.885 450.585 ;
  END
 END o117
 PIN o118
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 446.025 26.885 446.595 ;
  END
 END o118
 PIN o119
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 441.845 26.885 442.415 ;
  END
 END o119
 PIN o120
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 437.855 26.885 438.425 ;
  END
 END o120
 PIN o121
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 433.675 26.885 434.245 ;
  END
 END o121
 PIN o122
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 429.685 26.885 430.255 ;
  END
 END o122
 PIN o123
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 425.505 26.885 426.075 ;
  END
 END o123
 PIN o124
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 720.385 26.885 720.955 ;
  END
 END o124
 PIN o125
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 421.515 26.885 422.085 ;
  END
 END o125
 PIN o126
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 417.335 26.885 417.905 ;
  END
 END o126
 PIN o127
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 413.345 26.885 413.915 ;
  END
 END o127
 PIN o128
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 409.165 26.885 409.735 ;
  END
 END o128
 PIN o129
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 405.175 26.885 405.745 ;
  END
 END o129
 PIN o130
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 400.995 26.885 401.565 ;
  END
 END o130
 PIN o131
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 397.005 26.885 397.575 ;
  END
 END o131
 PIN o132
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 392.825 26.885 393.395 ;
  END
 END o132
 PIN o133
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 388.835 26.885 389.405 ;
  END
 END o133
 PIN o134
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 384.655 26.885 385.225 ;
  END
 END o134
 PIN o135
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 716.395 26.885 716.965 ;
  END
 END o135
 PIN o136
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 356.535 26.885 357.105 ;
  END
 END o136
 PIN o137
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 352.355 26.885 352.925 ;
  END
 END o137
 PIN o138
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 348.365 26.885 348.935 ;
  END
 END o138
 PIN o139
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 344.185 26.885 344.755 ;
  END
 END o139
 PIN o140
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 340.195 26.885 340.765 ;
  END
 END o140
 PIN o141
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 336.015 26.885 336.585 ;
  END
 END o141
 PIN o142
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 332.025 26.885 332.595 ;
  END
 END o142
 PIN o143
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 327.845 26.885 328.415 ;
  END
 END o143
 PIN o144
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 323.855 26.885 324.425 ;
  END
 END o144
 PIN o145
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 319.675 26.885 320.245 ;
  END
 END o145
 PIN o146
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 712.215 26.885 712.785 ;
  END
 END o146
 PIN o147
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 315.685 26.885 316.255 ;
  END
 END o147
 PIN o148
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 311.505 26.885 312.075 ;
  END
 END o148
 PIN o149
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 307.515 26.885 308.085 ;
  END
 END o149
 PIN o150
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 303.335 26.885 303.905 ;
  END
 END o150
 PIN o151
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 299.345 26.885 299.915 ;
  END
 END o151
 PIN o152
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 295.165 26.885 295.735 ;
  END
 END o152
 PIN o153
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 291.175 26.885 291.745 ;
  END
 END o153
 PIN o154
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 286.995 26.885 287.565 ;
  END
 END o154
 PIN o155
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 283.005 26.885 283.575 ;
  END
 END o155
 PIN o156
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 278.825 26.885 279.395 ;
  END
 END o156
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 381.805 3.705 382.375 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 364.705 3.705 365.275 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 376.485 3.705 377.055 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 381.425 4.465 381.995 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 382.185 4.465 382.755 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 382.565 3.705 383.135 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 372.875 3.705 373.445 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 359.765 3.705 360.335 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 365.465 3.705 366.035 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 363.375 3.705 363.945 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 360.905 3.705 361.475 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 359.385 4.465 359.955 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 13.015 382.945 13.585 383.515 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 13.015 369.645 13.585 370.215 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 750.785 26.885 751.355 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 746.605 26.885 747.175 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 709.935 26.885 710.505 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 254.885 26.885 255.455 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 250.705 26.885 251.275 ;
  END
 END i18
 PIN i19
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 246.715 26.885 247.285 ;
  END
 END i19
 PIN i20
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 242.535 26.885 243.105 ;
  END
 END i20
 PIN i21
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 238.545 26.885 239.115 ;
  END
 END i21
 PIN i22
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 234.365 26.885 234.935 ;
  END
 END i22
 PIN i23
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 230.375 26.885 230.945 ;
  END
 END i23
 PIN i24
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 226.195 26.885 226.765 ;
  END
 END i24
 PIN i25
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 222.205 26.885 222.775 ;
  END
 END i25
 PIN i26
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 218.025 26.885 218.595 ;
  END
 END i26
 PIN i27
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 705.755 26.885 706.325 ;
  END
 END i27
 PIN i28
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 214.035 26.885 214.605 ;
  END
 END i28
 PIN i29
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 209.855 26.885 210.425 ;
  END
 END i29
 PIN i30
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 205.865 26.885 206.435 ;
  END
 END i30
 PIN i31
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 201.685 26.885 202.255 ;
  END
 END i31
 PIN i32
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 197.695 26.885 198.265 ;
  END
 END i32
 PIN i33
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 193.515 26.885 194.085 ;
  END
 END i33
 PIN i34
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 189.525 26.885 190.095 ;
  END
 END i34
 PIN i35
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 185.345 26.885 185.915 ;
  END
 END i35
 PIN i36
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 181.355 26.885 181.925 ;
  END
 END i36
 PIN i37
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 172.045 26.885 172.615 ;
  END
 END i37
 PIN i38
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 701.765 26.885 702.335 ;
  END
 END i38
 PIN i39
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 168.055 26.885 168.625 ;
  END
 END i39
 PIN i40
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 163.875 26.885 164.445 ;
  END
 END i40
 PIN i41
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 159.885 26.885 160.455 ;
  END
 END i41
 PIN i42
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 155.705 26.885 156.275 ;
  END
 END i42
 PIN i43
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 151.715 26.885 152.285 ;
  END
 END i43
 PIN i44
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 147.535 26.885 148.105 ;
  END
 END i44
 PIN i45
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 143.545 26.885 144.115 ;
  END
 END i45
 PIN i46
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 139.365 26.885 139.935 ;
  END
 END i46
 PIN i47
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 135.375 26.885 135.945 ;
  END
 END i47
 PIN i48
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 131.195 26.885 131.765 ;
  END
 END i48
 PIN i49
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 697.585 26.885 698.155 ;
  END
 END i49
 PIN i50
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 127.205 26.885 127.775 ;
  END
 END i50
 PIN i51
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 123.025 26.885 123.595 ;
  END
 END i51
 PIN i52
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 119.035 26.885 119.605 ;
  END
 END i52
 PIN i53
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 114.855 26.885 115.425 ;
  END
 END i53
 PIN i54
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 110.865 26.885 111.435 ;
  END
 END i54
 PIN i55
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 106.685 26.885 107.255 ;
  END
 END i55
 PIN i56
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 102.695 26.885 103.265 ;
  END
 END i56
 PIN i57
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 98.515 26.885 99.085 ;
  END
 END i57
 PIN i58
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 76.285 26.885 76.855 ;
  END
 END i58
 PIN i59
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 72.105 26.885 72.675 ;
  END
 END i59
 PIN i60
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 693.595 26.885 694.165 ;
  END
 END i60
 PIN i61
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 68.115 26.885 68.685 ;
  END
 END i61
 PIN i62
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 63.935 26.885 64.505 ;
  END
 END i62
 PIN i63
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 59.945 26.885 60.515 ;
  END
 END i63
 PIN i64
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 55.765 26.885 56.335 ;
  END
 END i64
 PIN i65
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 51.775 26.885 52.345 ;
  END
 END i65
 PIN i66
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 47.595 26.885 48.165 ;
  END
 END i66
 PIN i67
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 43.605 26.885 44.175 ;
  END
 END i67
 PIN i68
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 39.425 26.885 39.995 ;
  END
 END i68
 PIN i69
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 35.435 26.885 36.005 ;
  END
 END i69
 PIN i70
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 31.255 26.885 31.825 ;
  END
 END i70
 PIN i71
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 689.415 26.885 689.985 ;
  END
 END i71
 PIN i72
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 27.265 26.885 27.835 ;
  END
 END i72
 PIN i73
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 23.085 26.885 23.655 ;
  END
 END i73
 PIN i74
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 19.095 26.885 19.665 ;
  END
 END i74
 PIN i75
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 14.915 26.885 15.485 ;
  END
 END i75
 PIN i76
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 10.925 26.885 11.495 ;
  END
 END i76
 PIN i77
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 6.745 26.885 7.315 ;
  END
 END i77
 PIN i78
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 2.755 26.885 3.325 ;
  END
 END i78
 PIN i79
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 685.425 26.885 685.995 ;
  END
 END i79
 PIN i80
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 681.245 26.885 681.815 ;
  END
 END i80
 PIN i81
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 677.255 26.885 677.825 ;
  END
 END i81
 PIN i82
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 673.075 26.885 673.645 ;
  END
 END i82
 PIN i83
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 742.615 26.885 743.185 ;
  END
 END i83
 PIN i84
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 650.845 26.885 651.415 ;
  END
 END i84
 PIN i85
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 646.665 26.885 647.235 ;
  END
 END i85
 PIN i86
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 642.675 26.885 643.245 ;
  END
 END i86
 PIN i87
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 638.495 26.885 639.065 ;
  END
 END i87
 PIN i88
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 634.505 26.885 635.075 ;
  END
 END i88
 PIN i89
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 630.325 26.885 630.895 ;
  END
 END i89
 PIN i90
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 626.335 26.885 626.905 ;
  END
 END i90
 PIN i91
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 622.155 26.885 622.725 ;
  END
 END i91
 PIN i92
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 618.165 26.885 618.735 ;
  END
 END i92
 PIN i93
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 613.985 26.885 614.555 ;
  END
 END i93
 PIN i94
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 738.435 26.885 739.005 ;
  END
 END i94
 PIN i95
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 609.995 26.885 610.565 ;
  END
 END i95
 PIN i96
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 605.815 26.885 606.385 ;
  END
 END i96
 PIN i97
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 601.825 26.885 602.395 ;
  END
 END i97
 PIN i98
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 597.645 26.885 598.215 ;
  END
 END i98
 PIN i99
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 593.655 26.885 594.225 ;
  END
 END i99
 PIN i100
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 589.475 26.885 590.045 ;
  END
 END i100
 PIN i101
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 585.485 26.885 586.055 ;
  END
 END i101
 PIN i102
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 581.305 26.885 581.875 ;
  END
 END i102
 PIN i103
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 577.315 26.885 577.885 ;
  END
 END i103
 PIN i104
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 573.135 26.885 573.705 ;
  END
 END i104
 PIN i105
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 734.445 26.885 735.015 ;
  END
 END i105
 PIN i106
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 564.015 26.885 564.585 ;
  END
 END i106
 PIN i107
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 559.835 26.885 560.405 ;
  END
 END i107
 PIN i108
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 555.845 26.885 556.415 ;
  END
 END i108
 PIN i109
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 551.665 26.885 552.235 ;
  END
 END i109
 PIN i110
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 547.675 26.885 548.245 ;
  END
 END i110
 PIN i111
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 543.495 26.885 544.065 ;
  END
 END i111
 PIN i112
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 539.505 26.885 540.075 ;
  END
 END i112
 PIN i113
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 535.325 26.885 535.895 ;
  END
 END i113
 PIN i114
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 531.335 26.885 531.905 ;
  END
 END i114
 PIN i115
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 527.155 26.885 527.725 ;
  END
 END i115
 PIN i116
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 730.265 26.885 730.835 ;
  END
 END i116
 PIN i117
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 523.165 26.885 523.735 ;
  END
 END i117
 PIN i118
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 518.985 26.885 519.555 ;
  END
 END i118
 PIN i119
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 514.995 26.885 515.565 ;
  END
 END i119
 PIN i120
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 510.815 26.885 511.385 ;
  END
 END i120
 PIN i121
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 506.825 26.885 507.395 ;
  END
 END i121
 PIN i122
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 502.645 26.885 503.215 ;
  END
 END i122
 PIN i123
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 498.655 26.885 499.225 ;
  END
 END i123
 PIN i124
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 494.475 26.885 495.045 ;
  END
 END i124
 PIN i125
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 490.485 26.885 491.055 ;
  END
 END i125
 PIN i126
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 486.305 26.885 486.875 ;
  END
 END i126
 PIN i127
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 726.275 26.885 726.845 ;
  END
 END i127
 PIN i128
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 464.075 26.885 464.645 ;
  END
 END i128
 PIN i129
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 459.895 26.885 460.465 ;
  END
 END i129
 PIN i130
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 455.905 26.885 456.475 ;
  END
 END i130
 PIN i131
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 451.725 26.885 452.295 ;
  END
 END i131
 PIN i132
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 447.735 26.885 448.305 ;
  END
 END i132
 PIN i133
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 443.555 26.885 444.125 ;
  END
 END i133
 PIN i134
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 439.565 26.885 440.135 ;
  END
 END i134
 PIN i135
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 435.385 26.885 435.955 ;
  END
 END i135
 PIN i136
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 431.395 26.885 431.965 ;
  END
 END i136
 PIN i137
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 427.215 26.885 427.785 ;
  END
 END i137
 PIN i138
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 722.095 26.885 722.665 ;
  END
 END i138
 PIN i139
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 423.225 26.885 423.795 ;
  END
 END i139
 PIN i140
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 419.045 26.885 419.615 ;
  END
 END i140
 PIN i141
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 415.055 26.885 415.625 ;
  END
 END i141
 PIN i142
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 410.875 26.885 411.445 ;
  END
 END i142
 PIN i143
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 406.885 26.885 407.455 ;
  END
 END i143
 PIN i144
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 402.705 26.885 403.275 ;
  END
 END i144
 PIN i145
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 398.715 26.885 399.285 ;
  END
 END i145
 PIN i146
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 394.535 26.885 395.105 ;
  END
 END i146
 PIN i147
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 390.545 26.885 391.115 ;
  END
 END i147
 PIN i148
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 386.365 26.885 386.935 ;
  END
 END i148
 PIN i149
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 718.105 26.885 718.675 ;
  END
 END i149
 PIN i150
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 354.825 26.885 355.395 ;
  END
 END i150
 PIN i151
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 350.645 26.885 351.215 ;
  END
 END i151
 PIN i152
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 346.655 26.885 347.225 ;
  END
 END i152
 PIN i153
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 342.475 26.885 343.045 ;
  END
 END i153
 PIN i154
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 338.485 26.885 339.055 ;
  END
 END i154
 PIN i155
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 334.305 26.885 334.875 ;
  END
 END i155
 PIN i156
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 330.315 26.885 330.885 ;
  END
 END i156
 PIN i157
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 326.135 26.885 326.705 ;
  END
 END i157
 PIN i158
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 322.145 26.885 322.715 ;
  END
 END i158
 PIN i159
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 317.965 26.885 318.535 ;
  END
 END i159
 PIN i160
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 713.925 26.885 714.495 ;
  END
 END i160
 PIN i161
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 313.975 26.885 314.545 ;
  END
 END i161
 PIN i162
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 309.795 26.885 310.365 ;
  END
 END i162
 PIN i163
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 305.805 26.885 306.375 ;
  END
 END i163
 PIN i164
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 301.625 26.885 302.195 ;
  END
 END i164
 PIN i165
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 297.635 26.885 298.205 ;
  END
 END i165
 PIN i166
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 293.455 26.885 294.025 ;
  END
 END i166
 PIN i167
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 289.465 26.885 290.035 ;
  END
 END i167
 PIN i168
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 285.285 26.885 285.855 ;
  END
 END i168
 PIN i169
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 281.295 26.885 281.865 ;
  END
 END i169
 PIN i170
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 277.115 26.885 277.685 ;
  END
 END i170
 PIN i171
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 695.305 27.645 695.875 ;
  END
 END i171
 PIN i172
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 691.315 27.645 691.885 ;
  END
 END i172
 PIN i173
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 687.135 27.645 687.705 ;
  END
 END i173
 PIN i174
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 707.655 27.645 708.225 ;
  END
 END i174
 PIN i175
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 703.475 27.645 704.045 ;
  END
 END i175
 PIN i176
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 628.045 27.645 628.615 ;
  END
 END i176
 PIN i177
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 624.055 27.645 624.625 ;
  END
 END i177
 PIN i178
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 619.875 27.645 620.445 ;
  END
 END i178
 PIN i179
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 615.885 27.645 616.455 ;
  END
 END i179
 PIN i180
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 611.705 27.645 612.275 ;
  END
 END i180
 PIN i181
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 508.535 27.645 509.105 ;
  END
 END i181
 PIN i182
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 504.545 27.645 505.115 ;
  END
 END i182
 PIN i183
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 500.365 27.645 500.935 ;
  END
 END i183
 PIN i184
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 520.885 27.645 521.455 ;
  END
 END i184
 PIN i185
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 516.705 27.645 517.275 ;
  END
 END i185
 PIN i186
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 441.275 27.645 441.845 ;
  END
 END i186
 PIN i187
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 437.285 27.645 437.855 ;
  END
 END i187
 PIN i188
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 433.105 27.645 433.675 ;
  END
 END i188
 PIN i189
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 429.115 27.645 429.685 ;
  END
 END i189
 PIN i190
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 424.935 27.645 425.505 ;
  END
 END i190
 PIN i191
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 299.915 27.645 300.485 ;
  END
 END i191
 PIN i192
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 303.905 27.645 304.475 ;
  END
 END i192
 PIN i193
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 308.085 27.645 308.655 ;
  END
 END i193
 PIN i194
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 312.075 27.645 312.645 ;
  END
 END i194
 PIN i195
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 316.255 27.645 316.825 ;
  END
 END i195
 PIN i196
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 232.655 27.645 233.225 ;
  END
 END i196
 PIN i197
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 236.645 27.645 237.215 ;
  END
 END i197
 PIN i198
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 240.825 27.645 241.395 ;
  END
 END i198
 PIN i199
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 220.305 27.645 220.875 ;
  END
 END i199
 PIN i200
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 224.485 27.645 225.055 ;
  END
 END i200
 PIN i201
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 121.315 27.645 121.885 ;
  END
 END i201
 PIN i202
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 125.305 27.645 125.875 ;
  END
 END i202
 PIN i203
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 129.485 27.645 130.055 ;
  END
 END i203
 PIN i204
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 133.475 27.645 134.045 ;
  END
 END i204
 PIN i205
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 137.655 27.645 138.225 ;
  END
 END i205
 PIN i206
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 54.055 27.645 54.625 ;
  END
 END i206
 PIN i207
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 58.045 27.645 58.615 ;
  END
 END i207
 PIN i208
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 62.225 27.645 62.795 ;
  END
 END i208
 PIN i209
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 41.705 27.645 42.275 ;
  END
 END i209
 PIN i210
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 45.885 27.645 46.455 ;
  END
 END i210
 PIN i211
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 699.485 27.645 700.055 ;
  END
 END i211
 PIN i212
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 632.225 27.645 632.795 ;
  END
 END i212
 PIN i213
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 512.715 27.645 513.285 ;
  END
 END i213
 PIN i214
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 445.455 27.645 446.025 ;
  END
 END i214
 PIN i215
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 295.735 27.645 296.305 ;
  END
 END i215
 PIN i216
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 228.475 27.645 229.045 ;
  END
 END i216
 PIN i217
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 117.135 27.645 117.705 ;
  END
 END i217
 PIN i218
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 49.875 27.645 50.445 ;
  END
 END i218
 PIN i219
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 17.955 382.945 18.525 383.515 ;
  END
 END i219
 PIN i220
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 17.955 369.645 18.525 370.215 ;
  END
 END i220
 PIN i221
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 750.215 27.645 750.785 ;
  END
 END i221
 PIN i222
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 746.035 27.645 746.605 ;
  END
 END i222
 PIN i223
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 709.365 27.645 709.935 ;
  END
 END i223
 PIN i224
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 255.455 27.645 256.025 ;
  END
 END i224
 PIN i225
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 251.275 27.645 251.845 ;
  END
 END i225
 PIN i226
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 247.285 27.645 247.855 ;
  END
 END i226
 PIN i227
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 243.105 27.645 243.675 ;
  END
 END i227
 PIN i228
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 239.115 27.645 239.685 ;
  END
 END i228
 PIN i229
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 234.935 27.645 235.505 ;
  END
 END i229
 PIN i230
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 230.945 27.645 231.515 ;
  END
 END i230
 PIN i231
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 226.765 27.645 227.335 ;
  END
 END i231
 PIN i232
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 222.775 27.645 223.345 ;
  END
 END i232
 PIN i233
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 218.595 27.645 219.165 ;
  END
 END i233
 PIN i234
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 705.185 27.645 705.755 ;
  END
 END i234
 PIN i235
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 214.605 27.645 215.175 ;
  END
 END i235
 PIN i236
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 210.425 27.645 210.995 ;
  END
 END i236
 PIN i237
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 206.435 27.645 207.005 ;
  END
 END i237
 PIN i238
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 202.255 27.645 202.825 ;
  END
 END i238
 PIN i239
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 198.265 27.645 198.835 ;
  END
 END i239
 PIN i240
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 194.085 27.645 194.655 ;
  END
 END i240
 PIN i241
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 190.095 27.645 190.665 ;
  END
 END i241
 PIN i242
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 185.915 27.645 186.485 ;
  END
 END i242
 PIN i243
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 181.925 27.645 182.495 ;
  END
 END i243
 PIN i244
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 172.615 27.645 173.185 ;
  END
 END i244
 PIN i245
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 701.195 27.645 701.765 ;
  END
 END i245
 PIN i246
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 168.625 27.645 169.195 ;
  END
 END i246
 PIN i247
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 164.445 27.645 165.015 ;
  END
 END i247
 PIN i248
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 160.455 27.645 161.025 ;
  END
 END i248
 PIN i249
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 156.275 27.645 156.845 ;
  END
 END i249
 PIN i250
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 152.285 27.645 152.855 ;
  END
 END i250
 PIN i251
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 148.105 27.645 148.675 ;
  END
 END i251
 PIN i252
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 144.115 27.645 144.685 ;
  END
 END i252
 PIN i253
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 139.935 27.645 140.505 ;
  END
 END i253
 PIN i254
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 135.945 27.645 136.515 ;
  END
 END i254
 PIN i255
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 131.765 27.645 132.335 ;
  END
 END i255
 PIN i256
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 697.015 27.645 697.585 ;
  END
 END i256
 PIN i257
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 127.775 27.645 128.345 ;
  END
 END i257
 PIN i258
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 123.595 27.645 124.165 ;
  END
 END i258
 PIN i259
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 119.605 27.645 120.175 ;
  END
 END i259
 PIN i260
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 115.425 27.645 115.995 ;
  END
 END i260
 PIN i261
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 111.435 27.645 112.005 ;
  END
 END i261
 PIN i262
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 107.255 27.645 107.825 ;
  END
 END i262
 PIN i263
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 103.265 27.645 103.835 ;
  END
 END i263
 PIN i264
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 99.085 27.645 99.655 ;
  END
 END i264
 PIN i265
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 76.855 27.645 77.425 ;
  END
 END i265
 PIN i266
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 72.675 27.645 73.245 ;
  END
 END i266
 PIN i267
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 693.025 27.645 693.595 ;
  END
 END i267
 PIN i268
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 68.685 27.645 69.255 ;
  END
 END i268
 PIN i269
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 64.505 27.645 65.075 ;
  END
 END i269
 PIN i270
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 60.515 27.645 61.085 ;
  END
 END i270
 PIN i271
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 56.335 27.645 56.905 ;
  END
 END i271
 PIN i272
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 52.345 27.645 52.915 ;
  END
 END i272
 PIN i273
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 48.165 27.645 48.735 ;
  END
 END i273
 PIN i274
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 44.175 27.645 44.745 ;
  END
 END i274
 PIN i275
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 39.995 27.645 40.565 ;
  END
 END i275
 PIN i276
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 36.005 27.645 36.575 ;
  END
 END i276
 PIN i277
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 31.825 27.645 32.395 ;
  END
 END i277
 PIN i278
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 688.845 27.645 689.415 ;
  END
 END i278
 PIN i279
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 27.835 27.645 28.405 ;
  END
 END i279
 PIN i280
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 23.655 27.645 24.225 ;
  END
 END i280
 PIN i281
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 19.665 27.645 20.235 ;
  END
 END i281
 PIN i282
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 15.485 27.645 16.055 ;
  END
 END i282
 PIN i283
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 11.495 27.645 12.065 ;
  END
 END i283
 PIN i284
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 7.315 27.645 7.885 ;
  END
 END i284
 PIN i285
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 3.325 27.645 3.895 ;
  END
 END i285
 PIN i286
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 684.855 27.645 685.425 ;
  END
 END i286
 PIN i287
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 680.675 27.645 681.245 ;
  END
 END i287
 PIN i288
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 676.685 27.645 677.255 ;
  END
 END i288
 PIN i289
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 672.505 27.645 673.075 ;
  END
 END i289
 PIN i290
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 742.045 27.645 742.615 ;
  END
 END i290
 PIN i291
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 650.275 27.645 650.845 ;
  END
 END i291
 PIN i292
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 646.095 27.645 646.665 ;
  END
 END i292
 PIN i293
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 642.105 27.645 642.675 ;
  END
 END i293
 PIN i294
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 637.925 27.645 638.495 ;
  END
 END i294
 PIN i295
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 633.935 27.645 634.505 ;
  END
 END i295
 PIN i296
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 629.755 27.645 630.325 ;
  END
 END i296
 PIN i297
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 625.765 27.645 626.335 ;
  END
 END i297
 PIN i298
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 621.585 27.645 622.155 ;
  END
 END i298
 PIN i299
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 617.595 27.645 618.165 ;
  END
 END i299
 PIN i300
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 613.415 27.645 613.985 ;
  END
 END i300
 PIN i301
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 737.865 27.645 738.435 ;
  END
 END i301
 PIN i302
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 609.425 27.645 609.995 ;
  END
 END i302
 PIN i303
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 605.245 27.645 605.815 ;
  END
 END i303
 PIN i304
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 601.255 27.645 601.825 ;
  END
 END i304
 PIN i305
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 597.075 27.645 597.645 ;
  END
 END i305
 PIN i306
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 593.085 27.645 593.655 ;
  END
 END i306
 PIN i307
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 588.905 27.645 589.475 ;
  END
 END i307
 PIN i308
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 584.915 27.645 585.485 ;
  END
 END i308
 PIN i309
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 580.735 27.645 581.305 ;
  END
 END i309
 PIN i310
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 576.745 27.645 577.315 ;
  END
 END i310
 PIN i311
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 572.565 27.645 573.135 ;
  END
 END i311
 PIN i312
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 733.875 27.645 734.445 ;
  END
 END i312
 PIN i313
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 563.445 27.645 564.015 ;
  END
 END i313
 PIN i314
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 559.265 27.645 559.835 ;
  END
 END i314
 PIN i315
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 555.275 27.645 555.845 ;
  END
 END i315
 PIN i316
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 551.095 27.645 551.665 ;
  END
 END i316
 PIN i317
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 547.105 27.645 547.675 ;
  END
 END i317
 PIN i318
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 542.925 27.645 543.495 ;
  END
 END i318
 PIN i319
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 538.935 27.645 539.505 ;
  END
 END i319
 PIN i320
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 534.755 27.645 535.325 ;
  END
 END i320
 PIN i321
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 530.765 27.645 531.335 ;
  END
 END i321
 PIN i322
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 526.585 27.645 527.155 ;
  END
 END i322
 PIN i323
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 729.695 27.645 730.265 ;
  END
 END i323
 PIN i324
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 522.595 27.645 523.165 ;
  END
 END i324
 PIN i325
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 518.415 27.645 518.985 ;
  END
 END i325
 PIN i326
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 514.425 27.645 514.995 ;
  END
 END i326
 PIN i327
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 510.245 27.645 510.815 ;
  END
 END i327
 PIN i328
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 506.255 27.645 506.825 ;
  END
 END i328
 PIN i329
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 502.075 27.645 502.645 ;
  END
 END i329
 PIN i330
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 498.085 27.645 498.655 ;
  END
 END i330
 PIN i331
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 493.905 27.645 494.475 ;
  END
 END i331
 PIN i332
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 489.915 27.645 490.485 ;
  END
 END i332
 PIN i333
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 485.735 27.645 486.305 ;
  END
 END i333
 PIN i334
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 725.705 27.645 726.275 ;
  END
 END i334
 PIN i335
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 463.505 27.645 464.075 ;
  END
 END i335
 PIN i336
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 459.325 27.645 459.895 ;
  END
 END i336
 PIN i337
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 455.335 27.645 455.905 ;
  END
 END i337
 PIN i338
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 451.155 27.645 451.725 ;
  END
 END i338
 PIN i339
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 447.165 27.645 447.735 ;
  END
 END i339
 PIN i340
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 442.985 27.645 443.555 ;
  END
 END i340
 PIN i341
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 438.995 27.645 439.565 ;
  END
 END i341
 PIN i342
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 434.815 27.645 435.385 ;
  END
 END i342
 PIN i343
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 430.825 27.645 431.395 ;
  END
 END i343
 PIN i344
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 426.645 27.645 427.215 ;
  END
 END i344
 PIN i345
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 721.525 27.645 722.095 ;
  END
 END i345
 PIN i346
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 422.655 27.645 423.225 ;
  END
 END i346
 PIN i347
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 418.475 27.645 419.045 ;
  END
 END i347
 PIN i348
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 414.485 27.645 415.055 ;
  END
 END i348
 PIN i349
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 410.305 27.645 410.875 ;
  END
 END i349
 PIN i350
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 406.315 27.645 406.885 ;
  END
 END i350
 PIN i351
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 402.135 27.645 402.705 ;
  END
 END i351
 PIN i352
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 398.145 27.645 398.715 ;
  END
 END i352
 PIN i353
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 393.965 27.645 394.535 ;
  END
 END i353
 PIN i354
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 389.975 27.645 390.545 ;
  END
 END i354
 PIN i355
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 385.795 27.645 386.365 ;
  END
 END i355
 PIN i356
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 717.535 27.645 718.105 ;
  END
 END i356
 PIN i357
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 355.395 27.645 355.965 ;
  END
 END i357
 PIN i358
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 351.215 27.645 351.785 ;
  END
 END i358
 PIN i359
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 347.225 27.645 347.795 ;
  END
 END i359
 PIN i360
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 343.045 27.645 343.615 ;
  END
 END i360
 PIN i361
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 339.055 27.645 339.625 ;
  END
 END i361
 PIN i362
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 334.875 27.645 335.445 ;
  END
 END i362
 PIN i363
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 330.885 27.645 331.455 ;
  END
 END i363
 PIN i364
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 326.705 27.645 327.275 ;
  END
 END i364
 PIN i365
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 322.715 27.645 323.285 ;
  END
 END i365
 PIN i366
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 318.535 27.645 319.105 ;
  END
 END i366
 PIN i367
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 713.355 27.645 713.925 ;
  END
 END i367
 PIN i368
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 314.545 27.645 315.115 ;
  END
 END i368
 PIN i369
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 310.365 27.645 310.935 ;
  END
 END i369
 PIN i370
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 306.375 27.645 306.945 ;
  END
 END i370
 PIN i371
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 302.195 27.645 302.765 ;
  END
 END i371
 PIN i372
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 298.205 27.645 298.775 ;
  END
 END i372
 PIN i373
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 294.025 27.645 294.595 ;
  END
 END i373
 PIN i374
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 290.035 27.645 290.605 ;
  END
 END i374
 PIN i375
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 285.855 27.645 286.425 ;
  END
 END i375
 PIN i376
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 281.865 27.645 282.435 ;
  END
 END i376
 PIN i377
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 277.685 27.645 278.255 ;
  END
 END i377
 PIN i378
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 375.345 3.705 375.915 ;
  END
 END i378
 PIN i379
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 374.965 4.465 375.535 ;
  END
 END i379
 PIN i380
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 749.645 28.405 750.215 ;
  END
 END i380
 PIN i381
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 745.465 28.405 746.035 ;
  END
 END i381
 PIN i382
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 708.795 28.405 709.365 ;
  END
 END i382
 PIN i383
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 256.025 28.405 256.595 ;
  END
 END i383
 PIN i384
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 251.845 28.405 252.415 ;
  END
 END i384
 PIN i385
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 247.855 28.405 248.425 ;
  END
 END i385
 PIN i386
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 243.675 28.405 244.245 ;
  END
 END i386
 PIN i387
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 239.685 28.405 240.255 ;
  END
 END i387
 PIN i388
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 235.505 28.405 236.075 ;
  END
 END i388
 PIN i389
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 231.515 28.405 232.085 ;
  END
 END i389
 PIN i390
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 227.335 28.405 227.905 ;
  END
 END i390
 PIN i391
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 223.345 28.405 223.915 ;
  END
 END i391
 PIN i392
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 219.165 28.405 219.735 ;
  END
 END i392
 PIN i393
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 704.615 28.405 705.185 ;
  END
 END i393
 PIN i394
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 215.175 28.405 215.745 ;
  END
 END i394
 PIN i395
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 210.995 28.405 211.565 ;
  END
 END i395
 PIN i396
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 207.005 28.405 207.575 ;
  END
 END i396
 PIN i397
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 202.825 28.405 203.395 ;
  END
 END i397
 PIN i398
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 198.835 28.405 199.405 ;
  END
 END i398
 PIN i399
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 194.655 28.405 195.225 ;
  END
 END i399
 PIN i400
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 190.665 28.405 191.235 ;
  END
 END i400
 PIN i401
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 186.485 28.405 187.055 ;
  END
 END i401
 PIN i402
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 182.495 28.405 183.065 ;
  END
 END i402
 PIN i403
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 173.185 28.405 173.755 ;
  END
 END i403
 PIN i404
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 700.625 28.405 701.195 ;
  END
 END i404
 PIN i405
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 169.195 28.405 169.765 ;
  END
 END i405
 PIN i406
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 165.015 28.405 165.585 ;
  END
 END i406
 PIN i407
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 161.025 28.405 161.595 ;
  END
 END i407
 PIN i408
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 156.845 28.405 157.415 ;
  END
 END i408
 PIN i409
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 152.855 28.405 153.425 ;
  END
 END i409
 PIN i410
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 148.675 28.405 149.245 ;
  END
 END i410
 PIN i411
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 144.685 28.405 145.255 ;
  END
 END i411
 PIN i412
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 140.505 28.405 141.075 ;
  END
 END i412
 PIN i413
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 136.515 28.405 137.085 ;
  END
 END i413
 PIN i414
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 132.335 28.405 132.905 ;
  END
 END i414
 PIN i415
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 696.445 28.405 697.015 ;
  END
 END i415
 PIN i416
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 128.345 28.405 128.915 ;
  END
 END i416
 PIN i417
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 124.165 28.405 124.735 ;
  END
 END i417
 PIN i418
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 120.175 28.405 120.745 ;
  END
 END i418
 PIN i419
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 115.995 28.405 116.565 ;
  END
 END i419
 PIN i420
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 112.005 28.405 112.575 ;
  END
 END i420
 PIN i421
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 107.825 28.405 108.395 ;
  END
 END i421
 PIN i422
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 103.835 28.405 104.405 ;
  END
 END i422
 PIN i423
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 99.655 28.405 100.225 ;
  END
 END i423
 PIN i424
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 77.425 28.405 77.995 ;
  END
 END i424
 PIN i425
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 73.245 28.405 73.815 ;
  END
 END i425
 PIN i426
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 692.455 28.405 693.025 ;
  END
 END i426
 PIN i427
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 69.255 28.405 69.825 ;
  END
 END i427
 PIN i428
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 65.075 28.405 65.645 ;
  END
 END i428
 PIN i429
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 61.085 28.405 61.655 ;
  END
 END i429
 PIN i430
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 56.905 28.405 57.475 ;
  END
 END i430
 PIN i431
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 52.915 28.405 53.485 ;
  END
 END i431
 PIN i432
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 48.735 28.405 49.305 ;
  END
 END i432
 PIN i433
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 44.745 28.405 45.315 ;
  END
 END i433
 PIN i434
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 40.565 28.405 41.135 ;
  END
 END i434
 PIN i435
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 36.575 28.405 37.145 ;
  END
 END i435
 PIN i436
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 32.395 28.405 32.965 ;
  END
 END i436
 PIN i437
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 688.275 28.405 688.845 ;
  END
 END i437
 PIN i438
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 28.405 28.405 28.975 ;
  END
 END i438
 PIN i439
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 24.225 28.405 24.795 ;
  END
 END i439
 PIN i440
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 20.235 28.405 20.805 ;
  END
 END i440
 PIN i441
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 16.055 28.405 16.625 ;
  END
 END i441
 PIN i442
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 12.065 28.405 12.635 ;
  END
 END i442
 PIN i443
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 7.885 28.405 8.455 ;
  END
 END i443
 PIN i444
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 3.895 28.405 4.465 ;
  END
 END i444
 PIN i445
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 684.285 28.405 684.855 ;
  END
 END i445
 PIN i446
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 680.105 28.405 680.675 ;
  END
 END i446
 PIN i447
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 676.115 28.405 676.685 ;
  END
 END i447
 PIN i448
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 671.935 28.405 672.505 ;
  END
 END i448
 PIN i449
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 741.475 28.405 742.045 ;
  END
 END i449
 PIN i450
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 649.705 28.405 650.275 ;
  END
 END i450
 PIN i451
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 645.525 28.405 646.095 ;
  END
 END i451
 PIN i452
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 641.535 28.405 642.105 ;
  END
 END i452
 PIN i453
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 637.355 28.405 637.925 ;
  END
 END i453
 PIN i454
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 633.365 28.405 633.935 ;
  END
 END i454
 PIN i455
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 629.185 28.405 629.755 ;
  END
 END i455
 PIN i456
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 625.195 28.405 625.765 ;
  END
 END i456
 PIN i457
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 621.015 28.405 621.585 ;
  END
 END i457
 PIN i458
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 617.025 28.405 617.595 ;
  END
 END i458
 PIN i459
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 612.845 28.405 613.415 ;
  END
 END i459
 PIN i460
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 737.295 28.405 737.865 ;
  END
 END i460
 PIN i461
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 608.855 28.405 609.425 ;
  END
 END i461
 PIN i462
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 604.675 28.405 605.245 ;
  END
 END i462
 PIN i463
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 600.685 28.405 601.255 ;
  END
 END i463
 PIN i464
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 596.505 28.405 597.075 ;
  END
 END i464
 PIN i465
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 592.515 28.405 593.085 ;
  END
 END i465
 PIN i466
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 588.335 28.405 588.905 ;
  END
 END i466
 PIN i467
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 584.345 28.405 584.915 ;
  END
 END i467
 PIN i468
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 580.165 28.405 580.735 ;
  END
 END i468
 PIN i469
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 576.175 28.405 576.745 ;
  END
 END i469
 PIN i470
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 571.995 28.405 572.565 ;
  END
 END i470
 PIN i471
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 733.305 28.405 733.875 ;
  END
 END i471
 PIN i472
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 562.875 28.405 563.445 ;
  END
 END i472
 PIN i473
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 558.695 28.405 559.265 ;
  END
 END i473
 PIN i474
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 554.705 28.405 555.275 ;
  END
 END i474
 PIN i475
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 550.525 28.405 551.095 ;
  END
 END i475
 PIN i476
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 546.535 28.405 547.105 ;
  END
 END i476
 PIN i477
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 542.355 28.405 542.925 ;
  END
 END i477
 PIN i478
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 538.365 28.405 538.935 ;
  END
 END i478
 PIN i479
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 534.185 28.405 534.755 ;
  END
 END i479
 PIN i480
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 530.195 28.405 530.765 ;
  END
 END i480
 PIN i481
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 526.015 28.405 526.585 ;
  END
 END i481
 PIN i482
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 729.125 28.405 729.695 ;
  END
 END i482
 PIN i483
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 522.025 28.405 522.595 ;
  END
 END i483
 PIN i484
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 517.845 28.405 518.415 ;
  END
 END i484
 PIN i485
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 513.855 28.405 514.425 ;
  END
 END i485
 PIN i486
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 509.675 28.405 510.245 ;
  END
 END i486
 PIN i487
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 505.685 28.405 506.255 ;
  END
 END i487
 PIN i488
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 501.505 28.405 502.075 ;
  END
 END i488
 PIN i489
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 497.515 28.405 498.085 ;
  END
 END i489
 PIN i490
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 493.335 28.405 493.905 ;
  END
 END i490
 PIN i491
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 489.345 28.405 489.915 ;
  END
 END i491
 PIN i492
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 485.165 28.405 485.735 ;
  END
 END i492
 PIN i493
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 725.135 28.405 725.705 ;
  END
 END i493
 PIN i494
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 462.935 28.405 463.505 ;
  END
 END i494
 PIN i495
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 458.755 28.405 459.325 ;
  END
 END i495
 PIN i496
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 454.765 28.405 455.335 ;
  END
 END i496
 PIN i497
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 450.585 28.405 451.155 ;
  END
 END i497
 PIN i498
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 446.595 28.405 447.165 ;
  END
 END i498
 PIN i499
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 442.415 28.405 442.985 ;
  END
 END i499
 PIN i500
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 438.425 28.405 438.995 ;
  END
 END i500
 PIN i501
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 434.245 28.405 434.815 ;
  END
 END i501
 PIN i502
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 430.255 28.405 430.825 ;
  END
 END i502
 PIN i503
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 426.075 28.405 426.645 ;
  END
 END i503
 PIN i504
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 720.955 28.405 721.525 ;
  END
 END i504
 PIN i505
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 422.085 28.405 422.655 ;
  END
 END i505
 PIN i506
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 417.905 28.405 418.475 ;
  END
 END i506
 PIN i507
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 413.915 28.405 414.485 ;
  END
 END i507
 PIN i508
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 409.735 28.405 410.305 ;
  END
 END i508
 PIN i509
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 405.745 28.405 406.315 ;
  END
 END i509
 PIN i510
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 401.565 28.405 402.135 ;
  END
 END i510
 PIN i511
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 397.575 28.405 398.145 ;
  END
 END i511
 PIN i512
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 393.395 28.405 393.965 ;
  END
 END i512
 PIN i513
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 389.405 28.405 389.975 ;
  END
 END i513
 PIN i514
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 385.225 28.405 385.795 ;
  END
 END i514
 PIN i515
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 716.965 28.405 717.535 ;
  END
 END i515
 PIN i516
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 355.965 28.405 356.535 ;
  END
 END i516
 PIN i517
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 351.785 28.405 352.355 ;
  END
 END i517
 PIN i518
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 347.795 28.405 348.365 ;
  END
 END i518
 PIN i519
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 343.615 28.405 344.185 ;
  END
 END i519
 PIN i520
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 339.625 28.405 340.195 ;
  END
 END i520
 PIN i521
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 335.445 28.405 336.015 ;
  END
 END i521
 PIN i522
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 331.455 28.405 332.025 ;
  END
 END i522
 PIN i523
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 327.275 28.405 327.845 ;
  END
 END i523
 PIN i524
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 323.285 28.405 323.855 ;
  END
 END i524
 PIN i525
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 319.105 28.405 319.675 ;
  END
 END i525
 PIN i526
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 712.785 28.405 713.355 ;
  END
 END i526
 PIN i527
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 315.115 28.405 315.685 ;
  END
 END i527
 PIN i528
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 310.935 28.405 311.505 ;
  END
 END i528
 PIN i529
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 306.945 28.405 307.515 ;
  END
 END i529
 PIN i530
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 302.765 28.405 303.335 ;
  END
 END i530
 PIN i531
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 298.775 28.405 299.345 ;
  END
 END i531
 PIN i532
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 294.595 28.405 295.165 ;
  END
 END i532
 PIN i533
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 290.605 28.405 291.175 ;
  END
 END i533
 PIN i534
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 286.425 28.405 286.995 ;
  END
 END i534
 PIN i535
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 282.435 28.405 283.005 ;
  END
 END i535
 PIN i536
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 278.255 28.405 278.825 ;
  END
 END i536
 PIN i537
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 4.275 382.945 4.845 383.515 ;
  END
 END i537
 PIN i538
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 5.415 382.945 5.985 383.515 ;
  END
 END i538
 PIN i539
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 6.935 382.945 7.505 383.515 ;
  END
 END i539
 PIN i540
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 8.835 382.945 9.405 383.515 ;
  END
 END i540
 PIN i541
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 4.275 369.645 4.845 370.215 ;
  END
 END i541
 PIN i542
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 5.415 369.645 5.985 370.215 ;
  END
 END i542
 PIN i543
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 6.935 369.645 7.505 370.215 ;
  END
 END i543
 PIN i544
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 8.835 369.645 9.405 370.215 ;
  END
 END i544
 OBS
  LAYER metal1 ;
   RECT 23.18 0.0 157.32 1.71 ;
   RECT 23.18 1.71 157.32 3.42 ;
   RECT 23.18 3.42 157.32 5.13 ;
   RECT 23.18 5.13 157.32 6.84 ;
   RECT 23.18 6.84 157.32 8.55 ;
   RECT 23.18 8.55 157.32 10.26 ;
   RECT 23.18 10.26 157.32 11.97 ;
   RECT 23.18 11.97 157.32 13.68 ;
   RECT 23.18 13.68 157.32 15.39 ;
   RECT 23.18 15.39 157.32 17.1 ;
   RECT 23.18 17.1 157.32 18.81 ;
   RECT 23.18 18.81 157.32 20.52 ;
   RECT 23.18 20.52 157.32 22.23 ;
   RECT 23.18 22.23 157.32 23.94 ;
   RECT 23.18 23.94 157.32 25.65 ;
   RECT 23.18 25.65 157.32 27.36 ;
   RECT 23.18 27.36 157.32 29.07 ;
   RECT 23.18 29.07 157.32 30.78 ;
   RECT 23.18 30.78 157.32 32.49 ;
   RECT 23.18 32.49 157.32 34.2 ;
   RECT 23.18 34.2 157.32 35.91 ;
   RECT 23.18 35.91 157.32 37.62 ;
   RECT 23.18 37.62 157.32 39.33 ;
   RECT 23.18 39.33 157.32 41.04 ;
   RECT 23.18 41.04 157.32 42.75 ;
   RECT 23.18 42.75 157.32 44.46 ;
   RECT 23.18 44.46 157.32 46.17 ;
   RECT 23.18 46.17 157.32 47.88 ;
   RECT 23.18 47.88 157.32 49.59 ;
   RECT 23.18 49.59 157.32 51.3 ;
   RECT 23.18 51.3 157.32 53.01 ;
   RECT 23.18 53.01 157.32 54.72 ;
   RECT 23.18 54.72 157.32 56.43 ;
   RECT 23.18 56.43 157.32 58.14 ;
   RECT 23.18 58.14 157.32 59.85 ;
   RECT 23.18 59.85 157.32 61.56 ;
   RECT 23.18 61.56 157.32 63.27 ;
   RECT 23.18 63.27 157.32 64.98 ;
   RECT 23.18 64.98 157.32 66.69 ;
   RECT 23.18 66.69 157.32 68.4 ;
   RECT 23.18 68.4 157.32 70.11 ;
   RECT 23.18 70.11 157.32 71.82 ;
   RECT 23.18 71.82 157.32 73.53 ;
   RECT 23.18 73.53 157.32 75.24 ;
   RECT 23.18 75.24 157.32 76.95 ;
   RECT 23.18 76.95 157.32 78.66 ;
   RECT 23.18 78.66 157.32 80.37 ;
   RECT 23.18 80.37 157.32 82.08 ;
   RECT 23.18 82.08 157.32 83.79 ;
   RECT 23.18 83.79 157.32 85.5 ;
   RECT 23.18 85.5 157.32 87.21 ;
   RECT 23.18 87.21 157.32 88.92 ;
   RECT 23.18 88.92 157.32 90.63 ;
   RECT 23.18 90.63 157.32 92.34 ;
   RECT 23.18 92.34 157.32 94.05 ;
   RECT 23.18 94.05 157.32 95.76 ;
   RECT 23.18 95.76 157.32 97.47 ;
   RECT 23.18 97.47 157.32 99.18 ;
   RECT 23.18 99.18 157.32 100.89 ;
   RECT 23.18 100.89 157.32 102.6 ;
   RECT 23.18 102.6 157.32 104.31 ;
   RECT 23.18 104.31 157.32 106.02 ;
   RECT 23.18 106.02 157.32 107.73 ;
   RECT 23.18 107.73 157.32 109.44 ;
   RECT 23.18 109.44 157.32 111.15 ;
   RECT 23.18 111.15 157.32 112.86 ;
   RECT 23.18 112.86 157.32 114.57 ;
   RECT 23.18 114.57 157.32 116.28 ;
   RECT 23.18 116.28 157.32 117.99 ;
   RECT 23.18 117.99 157.32 119.7 ;
   RECT 23.18 119.7 157.32 121.41 ;
   RECT 23.18 121.41 157.32 123.12 ;
   RECT 23.18 123.12 157.32 124.83 ;
   RECT 23.18 124.83 157.32 126.54 ;
   RECT 23.18 126.54 157.32 128.25 ;
   RECT 23.18 128.25 157.32 129.96 ;
   RECT 23.18 129.96 157.32 131.67 ;
   RECT 23.18 131.67 157.32 133.38 ;
   RECT 23.18 133.38 157.32 135.09 ;
   RECT 23.18 135.09 157.32 136.8 ;
   RECT 23.18 136.8 157.32 138.51 ;
   RECT 23.18 138.51 157.32 140.22 ;
   RECT 23.18 140.22 157.32 141.93 ;
   RECT 23.18 141.93 157.32 143.64 ;
   RECT 23.18 143.64 157.32 145.35 ;
   RECT 23.18 145.35 157.32 147.06 ;
   RECT 23.18 147.06 157.32 148.77 ;
   RECT 23.18 148.77 157.32 150.48 ;
   RECT 23.18 150.48 157.32 152.19 ;
   RECT 23.18 152.19 157.32 153.9 ;
   RECT 23.18 153.9 157.32 155.61 ;
   RECT 23.18 155.61 157.32 157.32 ;
   RECT 23.18 157.32 157.32 159.03 ;
   RECT 23.18 159.03 157.32 160.74 ;
   RECT 23.18 160.74 157.32 162.45 ;
   RECT 23.18 162.45 157.32 164.16 ;
   RECT 23.18 164.16 157.32 165.87 ;
   RECT 23.18 165.87 157.32 167.58 ;
   RECT 23.18 167.58 157.32 169.29 ;
   RECT 23.18 169.29 157.32 171.0 ;
   RECT 23.18 171.0 157.32 172.71 ;
   RECT 23.18 172.71 157.32 174.42 ;
   RECT 23.18 174.42 157.32 176.13 ;
   RECT 23.18 176.13 157.32 177.84 ;
   RECT 23.18 177.84 157.32 179.55 ;
   RECT 23.18 179.55 157.32 181.26 ;
   RECT 23.18 181.26 157.32 182.97 ;
   RECT 23.18 182.97 157.32 184.68 ;
   RECT 23.18 184.68 157.32 186.39 ;
   RECT 23.18 186.39 157.32 188.1 ;
   RECT 23.18 188.1 157.32 189.81 ;
   RECT 23.18 189.81 157.32 191.52 ;
   RECT 23.18 191.52 157.32 193.23 ;
   RECT 23.18 193.23 157.32 194.94 ;
   RECT 23.18 194.94 157.32 196.65 ;
   RECT 23.18 196.65 157.32 198.36 ;
   RECT 23.18 198.36 157.32 200.07 ;
   RECT 23.18 200.07 157.32 201.78 ;
   RECT 23.18 201.78 157.32 203.49 ;
   RECT 23.18 203.49 157.32 205.2 ;
   RECT 23.18 205.2 157.32 206.91 ;
   RECT 23.18 206.91 157.32 208.62 ;
   RECT 23.18 208.62 157.32 210.33 ;
   RECT 23.18 210.33 157.32 212.04 ;
   RECT 23.18 212.04 157.32 213.75 ;
   RECT 23.18 213.75 157.32 215.46 ;
   RECT 23.18 215.46 157.32 217.17 ;
   RECT 23.18 217.17 157.32 218.88 ;
   RECT 23.18 218.88 157.32 220.59 ;
   RECT 23.18 220.59 157.32 222.3 ;
   RECT 23.18 222.3 157.32 224.01 ;
   RECT 23.18 224.01 157.32 225.72 ;
   RECT 23.18 225.72 157.32 227.43 ;
   RECT 23.18 227.43 157.32 229.14 ;
   RECT 23.18 229.14 157.32 230.85 ;
   RECT 23.18 230.85 157.32 232.56 ;
   RECT 23.18 232.56 157.32 234.27 ;
   RECT 23.18 234.27 157.32 235.98 ;
   RECT 23.18 235.98 157.32 237.69 ;
   RECT 23.18 237.69 157.32 239.4 ;
   RECT 23.18 239.4 157.32 241.11 ;
   RECT 23.18 241.11 157.32 242.82 ;
   RECT 23.18 242.82 157.32 244.53 ;
   RECT 23.18 244.53 157.32 246.24 ;
   RECT 23.18 246.24 157.32 247.95 ;
   RECT 23.18 247.95 157.32 249.66 ;
   RECT 23.18 249.66 157.32 251.37 ;
   RECT 23.18 251.37 157.32 253.08 ;
   RECT 23.18 253.08 157.32 254.79 ;
   RECT 23.18 254.79 157.32 256.5 ;
   RECT 23.18 256.5 157.32 258.21 ;
   RECT 23.18 258.21 157.32 259.92 ;
   RECT 23.18 259.92 157.32 261.63 ;
   RECT 23.18 261.63 157.32 263.34 ;
   RECT 23.18 263.34 157.32 265.05 ;
   RECT 23.18 265.05 157.32 266.76 ;
   RECT 23.18 266.76 157.32 268.47 ;
   RECT 23.18 268.47 157.32 270.18 ;
   RECT 23.18 270.18 157.32 271.89 ;
   RECT 23.18 271.89 157.32 273.6 ;
   RECT 23.18 273.6 157.32 275.31 ;
   RECT 23.18 275.31 157.32 277.02 ;
   RECT 23.18 277.02 157.32 278.73 ;
   RECT 23.18 278.73 157.32 280.44 ;
   RECT 23.18 280.44 157.32 282.15 ;
   RECT 23.18 282.15 157.32 283.86 ;
   RECT 23.18 283.86 157.32 285.57 ;
   RECT 23.18 285.57 157.32 287.28 ;
   RECT 23.18 287.28 157.32 288.99 ;
   RECT 23.18 288.99 157.32 290.7 ;
   RECT 23.18 290.7 157.32 292.41 ;
   RECT 23.18 292.41 157.32 294.12 ;
   RECT 23.18 294.12 157.32 295.83 ;
   RECT 23.18 295.83 157.32 297.54 ;
   RECT 23.18 297.54 157.32 299.25 ;
   RECT 23.18 299.25 157.32 300.96 ;
   RECT 23.18 300.96 157.32 302.67 ;
   RECT 23.18 302.67 157.32 304.38 ;
   RECT 23.18 304.38 157.32 306.09 ;
   RECT 23.18 306.09 157.32 307.8 ;
   RECT 23.18 307.8 157.32 309.51 ;
   RECT 23.18 309.51 157.32 311.22 ;
   RECT 23.18 311.22 157.32 312.93 ;
   RECT 23.18 312.93 157.32 314.64 ;
   RECT 23.18 314.64 157.32 316.35 ;
   RECT 23.18 316.35 157.32 318.06 ;
   RECT 23.18 318.06 157.32 319.77 ;
   RECT 23.18 319.77 157.32 321.48 ;
   RECT 23.18 321.48 157.32 323.19 ;
   RECT 23.18 323.19 157.32 324.9 ;
   RECT 23.18 324.9 157.32 326.61 ;
   RECT 23.18 326.61 157.32 328.32 ;
   RECT 23.18 328.32 157.32 330.03 ;
   RECT 23.18 330.03 157.32 331.74 ;
   RECT 23.18 331.74 157.32 333.45 ;
   RECT 23.18 333.45 157.32 335.16 ;
   RECT 23.18 335.16 157.32 336.87 ;
   RECT 23.18 336.87 157.32 338.58 ;
   RECT 23.18 338.58 157.32 340.29 ;
   RECT 23.18 340.29 157.32 342.0 ;
   RECT 23.18 342.0 157.32 343.71 ;
   RECT 23.18 343.71 157.32 345.42 ;
   RECT 23.18 345.42 157.32 347.13 ;
   RECT 23.18 347.13 157.32 348.84 ;
   RECT 23.18 348.84 157.32 350.55 ;
   RECT 23.18 350.55 157.32 352.26 ;
   RECT 23.18 352.26 157.32 353.97 ;
   RECT 23.18 353.97 157.32 355.68 ;
   RECT 23.18 355.68 157.32 357.39 ;
   RECT 0.0 357.39 157.32 359.1 ;
   RECT 0.0 359.1 157.32 360.81 ;
   RECT 0.0 360.81 157.32 362.52 ;
   RECT 0.0 362.52 157.32 364.23 ;
   RECT 0.0 364.23 157.32 365.94 ;
   RECT 0.0 365.94 157.32 367.65 ;
   RECT 0.0 367.65 157.32 369.36 ;
   RECT 0.0 369.36 157.32 371.07 ;
   RECT 0.0 371.07 157.32 372.78 ;
   RECT 0.0 372.78 157.32 374.49 ;
   RECT 0.0 374.49 157.32 376.2 ;
   RECT 0.0 376.2 157.32 377.91 ;
   RECT 0.0 377.91 157.32 379.62 ;
   RECT 0.0 379.62 157.32 381.33 ;
   RECT 0.0 381.33 157.32 383.04 ;
   RECT 0.0 383.04 157.32 384.75 ;
   RECT 0.0 384.75 157.32 386.46 ;
   RECT 23.18 386.46 157.32 388.17 ;
   RECT 23.18 388.17 157.32 389.88 ;
   RECT 23.18 389.88 157.32 391.59 ;
   RECT 23.18 391.59 157.32 393.3 ;
   RECT 23.18 393.3 157.32 395.01 ;
   RECT 23.18 395.01 157.32 396.72 ;
   RECT 23.18 396.72 157.32 398.43 ;
   RECT 23.18 398.43 157.32 400.14 ;
   RECT 23.18 400.14 157.32 401.85 ;
   RECT 23.18 401.85 157.32 403.56 ;
   RECT 23.18 403.56 157.32 405.27 ;
   RECT 23.18 405.27 157.32 406.98 ;
   RECT 23.18 406.98 157.32 408.69 ;
   RECT 23.18 408.69 157.32 410.4 ;
   RECT 23.18 410.4 157.32 412.11 ;
   RECT 23.18 412.11 157.32 413.82 ;
   RECT 23.18 413.82 157.32 415.53 ;
   RECT 23.18 415.53 157.32 417.24 ;
   RECT 23.18 417.24 157.32 418.95 ;
   RECT 23.18 418.95 157.32 420.66 ;
   RECT 23.18 420.66 157.32 422.37 ;
   RECT 23.18 422.37 157.32 424.08 ;
   RECT 23.18 424.08 157.32 425.79 ;
   RECT 23.18 425.79 157.32 427.5 ;
   RECT 23.18 427.5 157.32 429.21 ;
   RECT 23.18 429.21 157.32 430.92 ;
   RECT 23.18 430.92 157.32 432.63 ;
   RECT 23.18 432.63 157.32 434.34 ;
   RECT 23.18 434.34 157.32 436.05 ;
   RECT 23.18 436.05 157.32 437.76 ;
   RECT 23.18 437.76 157.32 439.47 ;
   RECT 23.18 439.47 157.32 441.18 ;
   RECT 23.18 441.18 157.32 442.89 ;
   RECT 23.18 442.89 157.32 444.6 ;
   RECT 23.18 444.6 157.32 446.31 ;
   RECT 23.18 446.31 157.32 448.02 ;
   RECT 23.18 448.02 157.32 449.73 ;
   RECT 23.18 449.73 157.32 451.44 ;
   RECT 23.18 451.44 157.32 453.15 ;
   RECT 23.18 453.15 157.32 454.86 ;
   RECT 23.18 454.86 157.32 456.57 ;
   RECT 23.18 456.57 157.32 458.28 ;
   RECT 23.18 458.28 157.32 459.99 ;
   RECT 23.18 459.99 157.32 461.7 ;
   RECT 23.18 461.7 157.32 463.41 ;
   RECT 23.18 463.41 157.32 465.12 ;
   RECT 23.18 465.12 157.32 466.83 ;
   RECT 23.18 466.83 157.32 468.54 ;
   RECT 23.18 468.54 157.32 470.25 ;
   RECT 23.18 470.25 157.32 471.96 ;
   RECT 23.18 471.96 157.32 473.67 ;
   RECT 23.18 473.67 157.32 475.38 ;
   RECT 23.18 475.38 157.32 477.09 ;
   RECT 23.18 477.09 157.32 478.8 ;
   RECT 23.18 478.8 157.32 480.51 ;
   RECT 23.18 480.51 157.32 482.22 ;
   RECT 23.18 482.22 157.32 483.93 ;
   RECT 23.18 483.93 157.32 485.64 ;
   RECT 23.18 485.64 157.32 487.35 ;
   RECT 23.18 487.35 157.32 489.06 ;
   RECT 23.18 489.06 157.32 490.77 ;
   RECT 23.18 490.77 157.32 492.48 ;
   RECT 23.18 492.48 157.32 494.19 ;
   RECT 23.18 494.19 157.32 495.9 ;
   RECT 23.18 495.9 157.32 497.61 ;
   RECT 23.18 497.61 157.32 499.32 ;
   RECT 23.18 499.32 157.32 501.03 ;
   RECT 23.18 501.03 157.32 502.74 ;
   RECT 23.18 502.74 157.32 504.45 ;
   RECT 23.18 504.45 157.32 506.16 ;
   RECT 23.18 506.16 157.32 507.87 ;
   RECT 23.18 507.87 157.32 509.58 ;
   RECT 23.18 509.58 157.32 511.29 ;
   RECT 23.18 511.29 157.32 513.0 ;
   RECT 23.18 513.0 157.32 514.71 ;
   RECT 23.18 514.71 157.32 516.42 ;
   RECT 23.18 516.42 157.32 518.13 ;
   RECT 23.18 518.13 157.32 519.84 ;
   RECT 23.18 519.84 157.32 521.55 ;
   RECT 23.18 521.55 157.32 523.26 ;
   RECT 23.18 523.26 157.32 524.97 ;
   RECT 23.18 524.97 157.32 526.68 ;
   RECT 23.18 526.68 157.32 528.39 ;
   RECT 23.18 528.39 157.32 530.1 ;
   RECT 23.18 530.1 157.32 531.81 ;
   RECT 23.18 531.81 157.32 533.52 ;
   RECT 23.18 533.52 157.32 535.23 ;
   RECT 23.18 535.23 157.32 536.94 ;
   RECT 23.18 536.94 157.32 538.65 ;
   RECT 23.18 538.65 157.32 540.36 ;
   RECT 23.18 540.36 157.32 542.07 ;
   RECT 23.18 542.07 157.32 543.78 ;
   RECT 23.18 543.78 157.32 545.49 ;
   RECT 23.18 545.49 157.32 547.2 ;
   RECT 23.18 547.2 157.32 548.91 ;
   RECT 23.18 548.91 157.32 550.62 ;
   RECT 23.18 550.62 157.32 552.33 ;
   RECT 23.18 552.33 157.32 554.04 ;
   RECT 23.18 554.04 157.32 555.75 ;
   RECT 23.18 555.75 157.32 557.46 ;
   RECT 23.18 557.46 157.32 559.17 ;
   RECT 23.18 559.17 157.32 560.88 ;
   RECT 23.18 560.88 157.32 562.59 ;
   RECT 23.18 562.59 157.32 564.3 ;
   RECT 23.18 564.3 157.32 566.01 ;
   RECT 23.18 566.01 157.32 567.72 ;
   RECT 23.18 567.72 157.32 569.43 ;
   RECT 23.18 569.43 157.32 571.14 ;
   RECT 23.18 571.14 157.32 572.85 ;
   RECT 23.18 572.85 157.32 574.56 ;
   RECT 23.18 574.56 157.32 576.27 ;
   RECT 23.18 576.27 157.32 577.98 ;
   RECT 23.18 577.98 157.32 579.69 ;
   RECT 23.18 579.69 157.32 581.4 ;
   RECT 23.18 581.4 157.32 583.11 ;
   RECT 23.18 583.11 157.32 584.82 ;
   RECT 23.18 584.82 157.32 586.53 ;
   RECT 23.18 586.53 157.32 588.24 ;
   RECT 23.18 588.24 157.32 589.95 ;
   RECT 23.18 589.95 157.32 591.66 ;
   RECT 23.18 591.66 157.32 593.37 ;
   RECT 23.18 593.37 157.32 595.08 ;
   RECT 23.18 595.08 157.32 596.79 ;
   RECT 23.18 596.79 157.32 598.5 ;
   RECT 23.18 598.5 157.32 600.21 ;
   RECT 23.18 600.21 157.32 601.92 ;
   RECT 23.18 601.92 157.32 603.63 ;
   RECT 23.18 603.63 157.32 605.34 ;
   RECT 23.18 605.34 157.32 607.05 ;
   RECT 23.18 607.05 157.32 608.76 ;
   RECT 23.18 608.76 157.32 610.47 ;
   RECT 23.18 610.47 157.32 612.18 ;
   RECT 23.18 612.18 157.32 613.89 ;
   RECT 23.18 613.89 157.32 615.6 ;
   RECT 23.18 615.6 157.32 617.31 ;
   RECT 23.18 617.31 157.32 619.02 ;
   RECT 23.18 619.02 157.32 620.73 ;
   RECT 23.18 620.73 157.32 622.44 ;
   RECT 23.18 622.44 157.32 624.15 ;
   RECT 23.18 624.15 157.32 625.86 ;
   RECT 23.18 625.86 157.32 627.57 ;
   RECT 23.18 627.57 157.32 629.28 ;
   RECT 23.18 629.28 157.32 630.99 ;
   RECT 23.18 630.99 157.32 632.7 ;
   RECT 23.18 632.7 157.32 634.41 ;
   RECT 23.18 634.41 157.32 636.12 ;
   RECT 23.18 636.12 157.32 637.83 ;
   RECT 23.18 637.83 157.32 639.54 ;
   RECT 23.18 639.54 157.32 641.25 ;
   RECT 23.18 641.25 157.32 642.96 ;
   RECT 23.18 642.96 157.32 644.67 ;
   RECT 23.18 644.67 157.32 646.38 ;
   RECT 23.18 646.38 157.32 648.09 ;
   RECT 23.18 648.09 157.32 649.8 ;
   RECT 23.18 649.8 157.32 651.51 ;
   RECT 23.18 651.51 157.32 653.22 ;
   RECT 23.18 653.22 157.32 654.93 ;
   RECT 23.18 654.93 157.32 656.64 ;
   RECT 23.18 656.64 157.32 658.35 ;
   RECT 23.18 658.35 157.32 660.06 ;
   RECT 23.18 660.06 157.32 661.77 ;
   RECT 23.18 661.77 157.32 663.48 ;
   RECT 23.18 663.48 157.32 665.19 ;
   RECT 23.18 665.19 157.32 666.9 ;
   RECT 23.18 666.9 157.32 668.61 ;
   RECT 23.18 668.61 157.32 670.32 ;
   RECT 23.18 670.32 157.32 672.03 ;
   RECT 23.18 672.03 157.32 673.74 ;
   RECT 23.18 673.74 157.32 675.45 ;
   RECT 23.18 675.45 157.32 677.16 ;
   RECT 23.18 677.16 157.32 678.87 ;
   RECT 23.18 678.87 157.32 680.58 ;
   RECT 23.18 680.58 157.32 682.29 ;
   RECT 23.18 682.29 157.32 684.0 ;
   RECT 23.18 684.0 157.32 685.71 ;
   RECT 23.18 685.71 157.32 687.42 ;
   RECT 23.18 687.42 157.32 689.13 ;
   RECT 23.18 689.13 157.32 690.84 ;
   RECT 23.18 690.84 157.32 692.55 ;
   RECT 23.18 692.55 157.32 694.26 ;
   RECT 23.18 694.26 157.32 695.97 ;
   RECT 23.18 695.97 157.32 697.68 ;
   RECT 23.18 697.68 157.32 699.39 ;
   RECT 23.18 699.39 157.32 701.1 ;
   RECT 23.18 701.1 157.32 702.81 ;
   RECT 23.18 702.81 157.32 704.52 ;
   RECT 23.18 704.52 157.32 706.23 ;
   RECT 23.18 706.23 157.32 707.94 ;
   RECT 23.18 707.94 157.32 709.65 ;
   RECT 23.18 709.65 157.32 711.36 ;
   RECT 23.18 711.36 157.32 713.07 ;
   RECT 23.18 713.07 157.32 714.78 ;
   RECT 23.18 714.78 157.32 716.49 ;
   RECT 23.18 716.49 157.32 718.2 ;
   RECT 23.18 718.2 157.32 719.91 ;
   RECT 23.18 719.91 157.32 721.62 ;
   RECT 23.18 721.62 157.32 723.33 ;
   RECT 23.18 723.33 157.32 725.04 ;
   RECT 23.18 725.04 157.32 726.75 ;
   RECT 23.18 726.75 157.32 728.46 ;
   RECT 23.18 728.46 157.32 730.17 ;
   RECT 23.18 730.17 157.32 731.88 ;
   RECT 23.18 731.88 157.32 733.59 ;
   RECT 23.18 733.59 157.32 735.3 ;
   RECT 23.18 735.3 157.32 737.01 ;
   RECT 23.18 737.01 157.32 738.72 ;
   RECT 23.18 738.72 157.32 740.43 ;
   RECT 23.18 740.43 157.32 742.14 ;
   RECT 23.18 742.14 157.32 743.85 ;
   RECT 23.18 743.85 157.32 745.56 ;
   RECT 23.18 745.56 157.32 747.27 ;
   RECT 23.18 747.27 157.32 748.98 ;
   RECT 23.18 748.98 157.32 750.69 ;
   RECT 23.18 750.69 157.32 752.4 ;
   RECT 23.18 752.4 157.32 754.11 ;
   RECT 23.18 754.11 157.32 755.82 ;
  LAYER via1 ;
   RECT 23.18 0.0 157.32 1.71 ;
   RECT 23.18 1.71 157.32 3.42 ;
   RECT 23.18 3.42 157.32 5.13 ;
   RECT 23.18 5.13 157.32 6.84 ;
   RECT 23.18 6.84 157.32 8.55 ;
   RECT 23.18 8.55 157.32 10.26 ;
   RECT 23.18 10.26 157.32 11.97 ;
   RECT 23.18 11.97 157.32 13.68 ;
   RECT 23.18 13.68 157.32 15.39 ;
   RECT 23.18 15.39 157.32 17.1 ;
   RECT 23.18 17.1 157.32 18.81 ;
   RECT 23.18 18.81 157.32 20.52 ;
   RECT 23.18 20.52 157.32 22.23 ;
   RECT 23.18 22.23 157.32 23.94 ;
   RECT 23.18 23.94 157.32 25.65 ;
   RECT 23.18 25.65 157.32 27.36 ;
   RECT 23.18 27.36 157.32 29.07 ;
   RECT 23.18 29.07 157.32 30.78 ;
   RECT 23.18 30.78 157.32 32.49 ;
   RECT 23.18 32.49 157.32 34.2 ;
   RECT 23.18 34.2 157.32 35.91 ;
   RECT 23.18 35.91 157.32 37.62 ;
   RECT 23.18 37.62 157.32 39.33 ;
   RECT 23.18 39.33 157.32 41.04 ;
   RECT 23.18 41.04 157.32 42.75 ;
   RECT 23.18 42.75 157.32 44.46 ;
   RECT 23.18 44.46 157.32 46.17 ;
   RECT 23.18 46.17 157.32 47.88 ;
   RECT 23.18 47.88 157.32 49.59 ;
   RECT 23.18 49.59 157.32 51.3 ;
   RECT 23.18 51.3 157.32 53.01 ;
   RECT 23.18 53.01 157.32 54.72 ;
   RECT 23.18 54.72 157.32 56.43 ;
   RECT 23.18 56.43 157.32 58.14 ;
   RECT 23.18 58.14 157.32 59.85 ;
   RECT 23.18 59.85 157.32 61.56 ;
   RECT 23.18 61.56 157.32 63.27 ;
   RECT 23.18 63.27 157.32 64.98 ;
   RECT 23.18 64.98 157.32 66.69 ;
   RECT 23.18 66.69 157.32 68.4 ;
   RECT 23.18 68.4 157.32 70.11 ;
   RECT 23.18 70.11 157.32 71.82 ;
   RECT 23.18 71.82 157.32 73.53 ;
   RECT 23.18 73.53 157.32 75.24 ;
   RECT 23.18 75.24 157.32 76.95 ;
   RECT 23.18 76.95 157.32 78.66 ;
   RECT 23.18 78.66 157.32 80.37 ;
   RECT 23.18 80.37 157.32 82.08 ;
   RECT 23.18 82.08 157.32 83.79 ;
   RECT 23.18 83.79 157.32 85.5 ;
   RECT 23.18 85.5 157.32 87.21 ;
   RECT 23.18 87.21 157.32 88.92 ;
   RECT 23.18 88.92 157.32 90.63 ;
   RECT 23.18 90.63 157.32 92.34 ;
   RECT 23.18 92.34 157.32 94.05 ;
   RECT 23.18 94.05 157.32 95.76 ;
   RECT 23.18 95.76 157.32 97.47 ;
   RECT 23.18 97.47 157.32 99.18 ;
   RECT 23.18 99.18 157.32 100.89 ;
   RECT 23.18 100.89 157.32 102.6 ;
   RECT 23.18 102.6 157.32 104.31 ;
   RECT 23.18 104.31 157.32 106.02 ;
   RECT 23.18 106.02 157.32 107.73 ;
   RECT 23.18 107.73 157.32 109.44 ;
   RECT 23.18 109.44 157.32 111.15 ;
   RECT 23.18 111.15 157.32 112.86 ;
   RECT 23.18 112.86 157.32 114.57 ;
   RECT 23.18 114.57 157.32 116.28 ;
   RECT 23.18 116.28 157.32 117.99 ;
   RECT 23.18 117.99 157.32 119.7 ;
   RECT 23.18 119.7 157.32 121.41 ;
   RECT 23.18 121.41 157.32 123.12 ;
   RECT 23.18 123.12 157.32 124.83 ;
   RECT 23.18 124.83 157.32 126.54 ;
   RECT 23.18 126.54 157.32 128.25 ;
   RECT 23.18 128.25 157.32 129.96 ;
   RECT 23.18 129.96 157.32 131.67 ;
   RECT 23.18 131.67 157.32 133.38 ;
   RECT 23.18 133.38 157.32 135.09 ;
   RECT 23.18 135.09 157.32 136.8 ;
   RECT 23.18 136.8 157.32 138.51 ;
   RECT 23.18 138.51 157.32 140.22 ;
   RECT 23.18 140.22 157.32 141.93 ;
   RECT 23.18 141.93 157.32 143.64 ;
   RECT 23.18 143.64 157.32 145.35 ;
   RECT 23.18 145.35 157.32 147.06 ;
   RECT 23.18 147.06 157.32 148.77 ;
   RECT 23.18 148.77 157.32 150.48 ;
   RECT 23.18 150.48 157.32 152.19 ;
   RECT 23.18 152.19 157.32 153.9 ;
   RECT 23.18 153.9 157.32 155.61 ;
   RECT 23.18 155.61 157.32 157.32 ;
   RECT 23.18 157.32 157.32 159.03 ;
   RECT 23.18 159.03 157.32 160.74 ;
   RECT 23.18 160.74 157.32 162.45 ;
   RECT 23.18 162.45 157.32 164.16 ;
   RECT 23.18 164.16 157.32 165.87 ;
   RECT 23.18 165.87 157.32 167.58 ;
   RECT 23.18 167.58 157.32 169.29 ;
   RECT 23.18 169.29 157.32 171.0 ;
   RECT 23.18 171.0 157.32 172.71 ;
   RECT 23.18 172.71 157.32 174.42 ;
   RECT 23.18 174.42 157.32 176.13 ;
   RECT 23.18 176.13 157.32 177.84 ;
   RECT 23.18 177.84 157.32 179.55 ;
   RECT 23.18 179.55 157.32 181.26 ;
   RECT 23.18 181.26 157.32 182.97 ;
   RECT 23.18 182.97 157.32 184.68 ;
   RECT 23.18 184.68 157.32 186.39 ;
   RECT 23.18 186.39 157.32 188.1 ;
   RECT 23.18 188.1 157.32 189.81 ;
   RECT 23.18 189.81 157.32 191.52 ;
   RECT 23.18 191.52 157.32 193.23 ;
   RECT 23.18 193.23 157.32 194.94 ;
   RECT 23.18 194.94 157.32 196.65 ;
   RECT 23.18 196.65 157.32 198.36 ;
   RECT 23.18 198.36 157.32 200.07 ;
   RECT 23.18 200.07 157.32 201.78 ;
   RECT 23.18 201.78 157.32 203.49 ;
   RECT 23.18 203.49 157.32 205.2 ;
   RECT 23.18 205.2 157.32 206.91 ;
   RECT 23.18 206.91 157.32 208.62 ;
   RECT 23.18 208.62 157.32 210.33 ;
   RECT 23.18 210.33 157.32 212.04 ;
   RECT 23.18 212.04 157.32 213.75 ;
   RECT 23.18 213.75 157.32 215.46 ;
   RECT 23.18 215.46 157.32 217.17 ;
   RECT 23.18 217.17 157.32 218.88 ;
   RECT 23.18 218.88 157.32 220.59 ;
   RECT 23.18 220.59 157.32 222.3 ;
   RECT 23.18 222.3 157.32 224.01 ;
   RECT 23.18 224.01 157.32 225.72 ;
   RECT 23.18 225.72 157.32 227.43 ;
   RECT 23.18 227.43 157.32 229.14 ;
   RECT 23.18 229.14 157.32 230.85 ;
   RECT 23.18 230.85 157.32 232.56 ;
   RECT 23.18 232.56 157.32 234.27 ;
   RECT 23.18 234.27 157.32 235.98 ;
   RECT 23.18 235.98 157.32 237.69 ;
   RECT 23.18 237.69 157.32 239.4 ;
   RECT 23.18 239.4 157.32 241.11 ;
   RECT 23.18 241.11 157.32 242.82 ;
   RECT 23.18 242.82 157.32 244.53 ;
   RECT 23.18 244.53 157.32 246.24 ;
   RECT 23.18 246.24 157.32 247.95 ;
   RECT 23.18 247.95 157.32 249.66 ;
   RECT 23.18 249.66 157.32 251.37 ;
   RECT 23.18 251.37 157.32 253.08 ;
   RECT 23.18 253.08 157.32 254.79 ;
   RECT 23.18 254.79 157.32 256.5 ;
   RECT 23.18 256.5 157.32 258.21 ;
   RECT 23.18 258.21 157.32 259.92 ;
   RECT 23.18 259.92 157.32 261.63 ;
   RECT 23.18 261.63 157.32 263.34 ;
   RECT 23.18 263.34 157.32 265.05 ;
   RECT 23.18 265.05 157.32 266.76 ;
   RECT 23.18 266.76 157.32 268.47 ;
   RECT 23.18 268.47 157.32 270.18 ;
   RECT 23.18 270.18 157.32 271.89 ;
   RECT 23.18 271.89 157.32 273.6 ;
   RECT 23.18 273.6 157.32 275.31 ;
   RECT 23.18 275.31 157.32 277.02 ;
   RECT 23.18 277.02 157.32 278.73 ;
   RECT 23.18 278.73 157.32 280.44 ;
   RECT 23.18 280.44 157.32 282.15 ;
   RECT 23.18 282.15 157.32 283.86 ;
   RECT 23.18 283.86 157.32 285.57 ;
   RECT 23.18 285.57 157.32 287.28 ;
   RECT 23.18 287.28 157.32 288.99 ;
   RECT 23.18 288.99 157.32 290.7 ;
   RECT 23.18 290.7 157.32 292.41 ;
   RECT 23.18 292.41 157.32 294.12 ;
   RECT 23.18 294.12 157.32 295.83 ;
   RECT 23.18 295.83 157.32 297.54 ;
   RECT 23.18 297.54 157.32 299.25 ;
   RECT 23.18 299.25 157.32 300.96 ;
   RECT 23.18 300.96 157.32 302.67 ;
   RECT 23.18 302.67 157.32 304.38 ;
   RECT 23.18 304.38 157.32 306.09 ;
   RECT 23.18 306.09 157.32 307.8 ;
   RECT 23.18 307.8 157.32 309.51 ;
   RECT 23.18 309.51 157.32 311.22 ;
   RECT 23.18 311.22 157.32 312.93 ;
   RECT 23.18 312.93 157.32 314.64 ;
   RECT 23.18 314.64 157.32 316.35 ;
   RECT 23.18 316.35 157.32 318.06 ;
   RECT 23.18 318.06 157.32 319.77 ;
   RECT 23.18 319.77 157.32 321.48 ;
   RECT 23.18 321.48 157.32 323.19 ;
   RECT 23.18 323.19 157.32 324.9 ;
   RECT 23.18 324.9 157.32 326.61 ;
   RECT 23.18 326.61 157.32 328.32 ;
   RECT 23.18 328.32 157.32 330.03 ;
   RECT 23.18 330.03 157.32 331.74 ;
   RECT 23.18 331.74 157.32 333.45 ;
   RECT 23.18 333.45 157.32 335.16 ;
   RECT 23.18 335.16 157.32 336.87 ;
   RECT 23.18 336.87 157.32 338.58 ;
   RECT 23.18 338.58 157.32 340.29 ;
   RECT 23.18 340.29 157.32 342.0 ;
   RECT 23.18 342.0 157.32 343.71 ;
   RECT 23.18 343.71 157.32 345.42 ;
   RECT 23.18 345.42 157.32 347.13 ;
   RECT 23.18 347.13 157.32 348.84 ;
   RECT 23.18 348.84 157.32 350.55 ;
   RECT 23.18 350.55 157.32 352.26 ;
   RECT 23.18 352.26 157.32 353.97 ;
   RECT 23.18 353.97 157.32 355.68 ;
   RECT 23.18 355.68 157.32 357.39 ;
   RECT 0.0 357.39 157.32 359.1 ;
   RECT 0.0 359.1 157.32 360.81 ;
   RECT 0.0 360.81 157.32 362.52 ;
   RECT 0.0 362.52 157.32 364.23 ;
   RECT 0.0 364.23 157.32 365.94 ;
   RECT 0.0 365.94 157.32 367.65 ;
   RECT 0.0 367.65 157.32 369.36 ;
   RECT 0.0 369.36 157.32 371.07 ;
   RECT 0.0 371.07 157.32 372.78 ;
   RECT 0.0 372.78 157.32 374.49 ;
   RECT 0.0 374.49 157.32 376.2 ;
   RECT 0.0 376.2 157.32 377.91 ;
   RECT 0.0 377.91 157.32 379.62 ;
   RECT 0.0 379.62 157.32 381.33 ;
   RECT 0.0 381.33 157.32 383.04 ;
   RECT 0.0 383.04 157.32 384.75 ;
   RECT 0.0 384.75 157.32 386.46 ;
   RECT 23.18 386.46 157.32 388.17 ;
   RECT 23.18 388.17 157.32 389.88 ;
   RECT 23.18 389.88 157.32 391.59 ;
   RECT 23.18 391.59 157.32 393.3 ;
   RECT 23.18 393.3 157.32 395.01 ;
   RECT 23.18 395.01 157.32 396.72 ;
   RECT 23.18 396.72 157.32 398.43 ;
   RECT 23.18 398.43 157.32 400.14 ;
   RECT 23.18 400.14 157.32 401.85 ;
   RECT 23.18 401.85 157.32 403.56 ;
   RECT 23.18 403.56 157.32 405.27 ;
   RECT 23.18 405.27 157.32 406.98 ;
   RECT 23.18 406.98 157.32 408.69 ;
   RECT 23.18 408.69 157.32 410.4 ;
   RECT 23.18 410.4 157.32 412.11 ;
   RECT 23.18 412.11 157.32 413.82 ;
   RECT 23.18 413.82 157.32 415.53 ;
   RECT 23.18 415.53 157.32 417.24 ;
   RECT 23.18 417.24 157.32 418.95 ;
   RECT 23.18 418.95 157.32 420.66 ;
   RECT 23.18 420.66 157.32 422.37 ;
   RECT 23.18 422.37 157.32 424.08 ;
   RECT 23.18 424.08 157.32 425.79 ;
   RECT 23.18 425.79 157.32 427.5 ;
   RECT 23.18 427.5 157.32 429.21 ;
   RECT 23.18 429.21 157.32 430.92 ;
   RECT 23.18 430.92 157.32 432.63 ;
   RECT 23.18 432.63 157.32 434.34 ;
   RECT 23.18 434.34 157.32 436.05 ;
   RECT 23.18 436.05 157.32 437.76 ;
   RECT 23.18 437.76 157.32 439.47 ;
   RECT 23.18 439.47 157.32 441.18 ;
   RECT 23.18 441.18 157.32 442.89 ;
   RECT 23.18 442.89 157.32 444.6 ;
   RECT 23.18 444.6 157.32 446.31 ;
   RECT 23.18 446.31 157.32 448.02 ;
   RECT 23.18 448.02 157.32 449.73 ;
   RECT 23.18 449.73 157.32 451.44 ;
   RECT 23.18 451.44 157.32 453.15 ;
   RECT 23.18 453.15 157.32 454.86 ;
   RECT 23.18 454.86 157.32 456.57 ;
   RECT 23.18 456.57 157.32 458.28 ;
   RECT 23.18 458.28 157.32 459.99 ;
   RECT 23.18 459.99 157.32 461.7 ;
   RECT 23.18 461.7 157.32 463.41 ;
   RECT 23.18 463.41 157.32 465.12 ;
   RECT 23.18 465.12 157.32 466.83 ;
   RECT 23.18 466.83 157.32 468.54 ;
   RECT 23.18 468.54 157.32 470.25 ;
   RECT 23.18 470.25 157.32 471.96 ;
   RECT 23.18 471.96 157.32 473.67 ;
   RECT 23.18 473.67 157.32 475.38 ;
   RECT 23.18 475.38 157.32 477.09 ;
   RECT 23.18 477.09 157.32 478.8 ;
   RECT 23.18 478.8 157.32 480.51 ;
   RECT 23.18 480.51 157.32 482.22 ;
   RECT 23.18 482.22 157.32 483.93 ;
   RECT 23.18 483.93 157.32 485.64 ;
   RECT 23.18 485.64 157.32 487.35 ;
   RECT 23.18 487.35 157.32 489.06 ;
   RECT 23.18 489.06 157.32 490.77 ;
   RECT 23.18 490.77 157.32 492.48 ;
   RECT 23.18 492.48 157.32 494.19 ;
   RECT 23.18 494.19 157.32 495.9 ;
   RECT 23.18 495.9 157.32 497.61 ;
   RECT 23.18 497.61 157.32 499.32 ;
   RECT 23.18 499.32 157.32 501.03 ;
   RECT 23.18 501.03 157.32 502.74 ;
   RECT 23.18 502.74 157.32 504.45 ;
   RECT 23.18 504.45 157.32 506.16 ;
   RECT 23.18 506.16 157.32 507.87 ;
   RECT 23.18 507.87 157.32 509.58 ;
   RECT 23.18 509.58 157.32 511.29 ;
   RECT 23.18 511.29 157.32 513.0 ;
   RECT 23.18 513.0 157.32 514.71 ;
   RECT 23.18 514.71 157.32 516.42 ;
   RECT 23.18 516.42 157.32 518.13 ;
   RECT 23.18 518.13 157.32 519.84 ;
   RECT 23.18 519.84 157.32 521.55 ;
   RECT 23.18 521.55 157.32 523.26 ;
   RECT 23.18 523.26 157.32 524.97 ;
   RECT 23.18 524.97 157.32 526.68 ;
   RECT 23.18 526.68 157.32 528.39 ;
   RECT 23.18 528.39 157.32 530.1 ;
   RECT 23.18 530.1 157.32 531.81 ;
   RECT 23.18 531.81 157.32 533.52 ;
   RECT 23.18 533.52 157.32 535.23 ;
   RECT 23.18 535.23 157.32 536.94 ;
   RECT 23.18 536.94 157.32 538.65 ;
   RECT 23.18 538.65 157.32 540.36 ;
   RECT 23.18 540.36 157.32 542.07 ;
   RECT 23.18 542.07 157.32 543.78 ;
   RECT 23.18 543.78 157.32 545.49 ;
   RECT 23.18 545.49 157.32 547.2 ;
   RECT 23.18 547.2 157.32 548.91 ;
   RECT 23.18 548.91 157.32 550.62 ;
   RECT 23.18 550.62 157.32 552.33 ;
   RECT 23.18 552.33 157.32 554.04 ;
   RECT 23.18 554.04 157.32 555.75 ;
   RECT 23.18 555.75 157.32 557.46 ;
   RECT 23.18 557.46 157.32 559.17 ;
   RECT 23.18 559.17 157.32 560.88 ;
   RECT 23.18 560.88 157.32 562.59 ;
   RECT 23.18 562.59 157.32 564.3 ;
   RECT 23.18 564.3 157.32 566.01 ;
   RECT 23.18 566.01 157.32 567.72 ;
   RECT 23.18 567.72 157.32 569.43 ;
   RECT 23.18 569.43 157.32 571.14 ;
   RECT 23.18 571.14 157.32 572.85 ;
   RECT 23.18 572.85 157.32 574.56 ;
   RECT 23.18 574.56 157.32 576.27 ;
   RECT 23.18 576.27 157.32 577.98 ;
   RECT 23.18 577.98 157.32 579.69 ;
   RECT 23.18 579.69 157.32 581.4 ;
   RECT 23.18 581.4 157.32 583.11 ;
   RECT 23.18 583.11 157.32 584.82 ;
   RECT 23.18 584.82 157.32 586.53 ;
   RECT 23.18 586.53 157.32 588.24 ;
   RECT 23.18 588.24 157.32 589.95 ;
   RECT 23.18 589.95 157.32 591.66 ;
   RECT 23.18 591.66 157.32 593.37 ;
   RECT 23.18 593.37 157.32 595.08 ;
   RECT 23.18 595.08 157.32 596.79 ;
   RECT 23.18 596.79 157.32 598.5 ;
   RECT 23.18 598.5 157.32 600.21 ;
   RECT 23.18 600.21 157.32 601.92 ;
   RECT 23.18 601.92 157.32 603.63 ;
   RECT 23.18 603.63 157.32 605.34 ;
   RECT 23.18 605.34 157.32 607.05 ;
   RECT 23.18 607.05 157.32 608.76 ;
   RECT 23.18 608.76 157.32 610.47 ;
   RECT 23.18 610.47 157.32 612.18 ;
   RECT 23.18 612.18 157.32 613.89 ;
   RECT 23.18 613.89 157.32 615.6 ;
   RECT 23.18 615.6 157.32 617.31 ;
   RECT 23.18 617.31 157.32 619.02 ;
   RECT 23.18 619.02 157.32 620.73 ;
   RECT 23.18 620.73 157.32 622.44 ;
   RECT 23.18 622.44 157.32 624.15 ;
   RECT 23.18 624.15 157.32 625.86 ;
   RECT 23.18 625.86 157.32 627.57 ;
   RECT 23.18 627.57 157.32 629.28 ;
   RECT 23.18 629.28 157.32 630.99 ;
   RECT 23.18 630.99 157.32 632.7 ;
   RECT 23.18 632.7 157.32 634.41 ;
   RECT 23.18 634.41 157.32 636.12 ;
   RECT 23.18 636.12 157.32 637.83 ;
   RECT 23.18 637.83 157.32 639.54 ;
   RECT 23.18 639.54 157.32 641.25 ;
   RECT 23.18 641.25 157.32 642.96 ;
   RECT 23.18 642.96 157.32 644.67 ;
   RECT 23.18 644.67 157.32 646.38 ;
   RECT 23.18 646.38 157.32 648.09 ;
   RECT 23.18 648.09 157.32 649.8 ;
   RECT 23.18 649.8 157.32 651.51 ;
   RECT 23.18 651.51 157.32 653.22 ;
   RECT 23.18 653.22 157.32 654.93 ;
   RECT 23.18 654.93 157.32 656.64 ;
   RECT 23.18 656.64 157.32 658.35 ;
   RECT 23.18 658.35 157.32 660.06 ;
   RECT 23.18 660.06 157.32 661.77 ;
   RECT 23.18 661.77 157.32 663.48 ;
   RECT 23.18 663.48 157.32 665.19 ;
   RECT 23.18 665.19 157.32 666.9 ;
   RECT 23.18 666.9 157.32 668.61 ;
   RECT 23.18 668.61 157.32 670.32 ;
   RECT 23.18 670.32 157.32 672.03 ;
   RECT 23.18 672.03 157.32 673.74 ;
   RECT 23.18 673.74 157.32 675.45 ;
   RECT 23.18 675.45 157.32 677.16 ;
   RECT 23.18 677.16 157.32 678.87 ;
   RECT 23.18 678.87 157.32 680.58 ;
   RECT 23.18 680.58 157.32 682.29 ;
   RECT 23.18 682.29 157.32 684.0 ;
   RECT 23.18 684.0 157.32 685.71 ;
   RECT 23.18 685.71 157.32 687.42 ;
   RECT 23.18 687.42 157.32 689.13 ;
   RECT 23.18 689.13 157.32 690.84 ;
   RECT 23.18 690.84 157.32 692.55 ;
   RECT 23.18 692.55 157.32 694.26 ;
   RECT 23.18 694.26 157.32 695.97 ;
   RECT 23.18 695.97 157.32 697.68 ;
   RECT 23.18 697.68 157.32 699.39 ;
   RECT 23.18 699.39 157.32 701.1 ;
   RECT 23.18 701.1 157.32 702.81 ;
   RECT 23.18 702.81 157.32 704.52 ;
   RECT 23.18 704.52 157.32 706.23 ;
   RECT 23.18 706.23 157.32 707.94 ;
   RECT 23.18 707.94 157.32 709.65 ;
   RECT 23.18 709.65 157.32 711.36 ;
   RECT 23.18 711.36 157.32 713.07 ;
   RECT 23.18 713.07 157.32 714.78 ;
   RECT 23.18 714.78 157.32 716.49 ;
   RECT 23.18 716.49 157.32 718.2 ;
   RECT 23.18 718.2 157.32 719.91 ;
   RECT 23.18 719.91 157.32 721.62 ;
   RECT 23.18 721.62 157.32 723.33 ;
   RECT 23.18 723.33 157.32 725.04 ;
   RECT 23.18 725.04 157.32 726.75 ;
   RECT 23.18 726.75 157.32 728.46 ;
   RECT 23.18 728.46 157.32 730.17 ;
   RECT 23.18 730.17 157.32 731.88 ;
   RECT 23.18 731.88 157.32 733.59 ;
   RECT 23.18 733.59 157.32 735.3 ;
   RECT 23.18 735.3 157.32 737.01 ;
   RECT 23.18 737.01 157.32 738.72 ;
   RECT 23.18 738.72 157.32 740.43 ;
   RECT 23.18 740.43 157.32 742.14 ;
   RECT 23.18 742.14 157.32 743.85 ;
   RECT 23.18 743.85 157.32 745.56 ;
   RECT 23.18 745.56 157.32 747.27 ;
   RECT 23.18 747.27 157.32 748.98 ;
   RECT 23.18 748.98 157.32 750.69 ;
   RECT 23.18 750.69 157.32 752.4 ;
   RECT 23.18 752.4 157.32 754.11 ;
   RECT 23.18 754.11 157.32 755.82 ;
  LAYER metal2 ;
   RECT 23.18 0.0 157.32 1.71 ;
   RECT 23.18 1.71 157.32 3.42 ;
   RECT 23.18 3.42 157.32 5.13 ;
   RECT 23.18 5.13 157.32 6.84 ;
   RECT 23.18 6.84 157.32 8.55 ;
   RECT 23.18 8.55 157.32 10.26 ;
   RECT 23.18 10.26 157.32 11.97 ;
   RECT 23.18 11.97 157.32 13.68 ;
   RECT 23.18 13.68 157.32 15.39 ;
   RECT 23.18 15.39 157.32 17.1 ;
   RECT 23.18 17.1 157.32 18.81 ;
   RECT 23.18 18.81 157.32 20.52 ;
   RECT 23.18 20.52 157.32 22.23 ;
   RECT 23.18 22.23 157.32 23.94 ;
   RECT 23.18 23.94 157.32 25.65 ;
   RECT 23.18 25.65 157.32 27.36 ;
   RECT 23.18 27.36 157.32 29.07 ;
   RECT 23.18 29.07 157.32 30.78 ;
   RECT 23.18 30.78 157.32 32.49 ;
   RECT 23.18 32.49 157.32 34.2 ;
   RECT 23.18 34.2 157.32 35.91 ;
   RECT 23.18 35.91 157.32 37.62 ;
   RECT 23.18 37.62 157.32 39.33 ;
   RECT 23.18 39.33 157.32 41.04 ;
   RECT 23.18 41.04 157.32 42.75 ;
   RECT 23.18 42.75 157.32 44.46 ;
   RECT 23.18 44.46 157.32 46.17 ;
   RECT 23.18 46.17 157.32 47.88 ;
   RECT 23.18 47.88 157.32 49.59 ;
   RECT 23.18 49.59 157.32 51.3 ;
   RECT 23.18 51.3 157.32 53.01 ;
   RECT 23.18 53.01 157.32 54.72 ;
   RECT 23.18 54.72 157.32 56.43 ;
   RECT 23.18 56.43 157.32 58.14 ;
   RECT 23.18 58.14 157.32 59.85 ;
   RECT 23.18 59.85 157.32 61.56 ;
   RECT 23.18 61.56 157.32 63.27 ;
   RECT 23.18 63.27 157.32 64.98 ;
   RECT 23.18 64.98 157.32 66.69 ;
   RECT 23.18 66.69 157.32 68.4 ;
   RECT 23.18 68.4 157.32 70.11 ;
   RECT 23.18 70.11 157.32 71.82 ;
   RECT 23.18 71.82 157.32 73.53 ;
   RECT 23.18 73.53 157.32 75.24 ;
   RECT 23.18 75.24 157.32 76.95 ;
   RECT 23.18 76.95 157.32 78.66 ;
   RECT 23.18 78.66 157.32 80.37 ;
   RECT 23.18 80.37 157.32 82.08 ;
   RECT 23.18 82.08 157.32 83.79 ;
   RECT 23.18 83.79 157.32 85.5 ;
   RECT 23.18 85.5 157.32 87.21 ;
   RECT 23.18 87.21 157.32 88.92 ;
   RECT 23.18 88.92 157.32 90.63 ;
   RECT 23.18 90.63 157.32 92.34 ;
   RECT 23.18 92.34 157.32 94.05 ;
   RECT 23.18 94.05 157.32 95.76 ;
   RECT 23.18 95.76 157.32 97.47 ;
   RECT 23.18 97.47 157.32 99.18 ;
   RECT 23.18 99.18 157.32 100.89 ;
   RECT 23.18 100.89 157.32 102.6 ;
   RECT 23.18 102.6 157.32 104.31 ;
   RECT 23.18 104.31 157.32 106.02 ;
   RECT 23.18 106.02 157.32 107.73 ;
   RECT 23.18 107.73 157.32 109.44 ;
   RECT 23.18 109.44 157.32 111.15 ;
   RECT 23.18 111.15 157.32 112.86 ;
   RECT 23.18 112.86 157.32 114.57 ;
   RECT 23.18 114.57 157.32 116.28 ;
   RECT 23.18 116.28 157.32 117.99 ;
   RECT 23.18 117.99 157.32 119.7 ;
   RECT 23.18 119.7 157.32 121.41 ;
   RECT 23.18 121.41 157.32 123.12 ;
   RECT 23.18 123.12 157.32 124.83 ;
   RECT 23.18 124.83 157.32 126.54 ;
   RECT 23.18 126.54 157.32 128.25 ;
   RECT 23.18 128.25 157.32 129.96 ;
   RECT 23.18 129.96 157.32 131.67 ;
   RECT 23.18 131.67 157.32 133.38 ;
   RECT 23.18 133.38 157.32 135.09 ;
   RECT 23.18 135.09 157.32 136.8 ;
   RECT 23.18 136.8 157.32 138.51 ;
   RECT 23.18 138.51 157.32 140.22 ;
   RECT 23.18 140.22 157.32 141.93 ;
   RECT 23.18 141.93 157.32 143.64 ;
   RECT 23.18 143.64 157.32 145.35 ;
   RECT 23.18 145.35 157.32 147.06 ;
   RECT 23.18 147.06 157.32 148.77 ;
   RECT 23.18 148.77 157.32 150.48 ;
   RECT 23.18 150.48 157.32 152.19 ;
   RECT 23.18 152.19 157.32 153.9 ;
   RECT 23.18 153.9 157.32 155.61 ;
   RECT 23.18 155.61 157.32 157.32 ;
   RECT 23.18 157.32 157.32 159.03 ;
   RECT 23.18 159.03 157.32 160.74 ;
   RECT 23.18 160.74 157.32 162.45 ;
   RECT 23.18 162.45 157.32 164.16 ;
   RECT 23.18 164.16 157.32 165.87 ;
   RECT 23.18 165.87 157.32 167.58 ;
   RECT 23.18 167.58 157.32 169.29 ;
   RECT 23.18 169.29 157.32 171.0 ;
   RECT 23.18 171.0 157.32 172.71 ;
   RECT 23.18 172.71 157.32 174.42 ;
   RECT 23.18 174.42 157.32 176.13 ;
   RECT 23.18 176.13 157.32 177.84 ;
   RECT 23.18 177.84 157.32 179.55 ;
   RECT 23.18 179.55 157.32 181.26 ;
   RECT 23.18 181.26 157.32 182.97 ;
   RECT 23.18 182.97 157.32 184.68 ;
   RECT 23.18 184.68 157.32 186.39 ;
   RECT 23.18 186.39 157.32 188.1 ;
   RECT 23.18 188.1 157.32 189.81 ;
   RECT 23.18 189.81 157.32 191.52 ;
   RECT 23.18 191.52 157.32 193.23 ;
   RECT 23.18 193.23 157.32 194.94 ;
   RECT 23.18 194.94 157.32 196.65 ;
   RECT 23.18 196.65 157.32 198.36 ;
   RECT 23.18 198.36 157.32 200.07 ;
   RECT 23.18 200.07 157.32 201.78 ;
   RECT 23.18 201.78 157.32 203.49 ;
   RECT 23.18 203.49 157.32 205.2 ;
   RECT 23.18 205.2 157.32 206.91 ;
   RECT 23.18 206.91 157.32 208.62 ;
   RECT 23.18 208.62 157.32 210.33 ;
   RECT 23.18 210.33 157.32 212.04 ;
   RECT 23.18 212.04 157.32 213.75 ;
   RECT 23.18 213.75 157.32 215.46 ;
   RECT 23.18 215.46 157.32 217.17 ;
   RECT 23.18 217.17 157.32 218.88 ;
   RECT 23.18 218.88 157.32 220.59 ;
   RECT 23.18 220.59 157.32 222.3 ;
   RECT 23.18 222.3 157.32 224.01 ;
   RECT 23.18 224.01 157.32 225.72 ;
   RECT 23.18 225.72 157.32 227.43 ;
   RECT 23.18 227.43 157.32 229.14 ;
   RECT 23.18 229.14 157.32 230.85 ;
   RECT 23.18 230.85 157.32 232.56 ;
   RECT 23.18 232.56 157.32 234.27 ;
   RECT 23.18 234.27 157.32 235.98 ;
   RECT 23.18 235.98 157.32 237.69 ;
   RECT 23.18 237.69 157.32 239.4 ;
   RECT 23.18 239.4 157.32 241.11 ;
   RECT 23.18 241.11 157.32 242.82 ;
   RECT 23.18 242.82 157.32 244.53 ;
   RECT 23.18 244.53 157.32 246.24 ;
   RECT 23.18 246.24 157.32 247.95 ;
   RECT 23.18 247.95 157.32 249.66 ;
   RECT 23.18 249.66 157.32 251.37 ;
   RECT 23.18 251.37 157.32 253.08 ;
   RECT 23.18 253.08 157.32 254.79 ;
   RECT 23.18 254.79 157.32 256.5 ;
   RECT 23.18 256.5 157.32 258.21 ;
   RECT 23.18 258.21 157.32 259.92 ;
   RECT 23.18 259.92 157.32 261.63 ;
   RECT 23.18 261.63 157.32 263.34 ;
   RECT 23.18 263.34 157.32 265.05 ;
   RECT 23.18 265.05 157.32 266.76 ;
   RECT 23.18 266.76 157.32 268.47 ;
   RECT 23.18 268.47 157.32 270.18 ;
   RECT 23.18 270.18 157.32 271.89 ;
   RECT 23.18 271.89 157.32 273.6 ;
   RECT 23.18 273.6 157.32 275.31 ;
   RECT 23.18 275.31 157.32 277.02 ;
   RECT 23.18 277.02 157.32 278.73 ;
   RECT 23.18 278.73 157.32 280.44 ;
   RECT 23.18 280.44 157.32 282.15 ;
   RECT 23.18 282.15 157.32 283.86 ;
   RECT 23.18 283.86 157.32 285.57 ;
   RECT 23.18 285.57 157.32 287.28 ;
   RECT 23.18 287.28 157.32 288.99 ;
   RECT 23.18 288.99 157.32 290.7 ;
   RECT 23.18 290.7 157.32 292.41 ;
   RECT 23.18 292.41 157.32 294.12 ;
   RECT 23.18 294.12 157.32 295.83 ;
   RECT 23.18 295.83 157.32 297.54 ;
   RECT 23.18 297.54 157.32 299.25 ;
   RECT 23.18 299.25 157.32 300.96 ;
   RECT 23.18 300.96 157.32 302.67 ;
   RECT 23.18 302.67 157.32 304.38 ;
   RECT 23.18 304.38 157.32 306.09 ;
   RECT 23.18 306.09 157.32 307.8 ;
   RECT 23.18 307.8 157.32 309.51 ;
   RECT 23.18 309.51 157.32 311.22 ;
   RECT 23.18 311.22 157.32 312.93 ;
   RECT 23.18 312.93 157.32 314.64 ;
   RECT 23.18 314.64 157.32 316.35 ;
   RECT 23.18 316.35 157.32 318.06 ;
   RECT 23.18 318.06 157.32 319.77 ;
   RECT 23.18 319.77 157.32 321.48 ;
   RECT 23.18 321.48 157.32 323.19 ;
   RECT 23.18 323.19 157.32 324.9 ;
   RECT 23.18 324.9 157.32 326.61 ;
   RECT 23.18 326.61 157.32 328.32 ;
   RECT 23.18 328.32 157.32 330.03 ;
   RECT 23.18 330.03 157.32 331.74 ;
   RECT 23.18 331.74 157.32 333.45 ;
   RECT 23.18 333.45 157.32 335.16 ;
   RECT 23.18 335.16 157.32 336.87 ;
   RECT 23.18 336.87 157.32 338.58 ;
   RECT 23.18 338.58 157.32 340.29 ;
   RECT 23.18 340.29 157.32 342.0 ;
   RECT 23.18 342.0 157.32 343.71 ;
   RECT 23.18 343.71 157.32 345.42 ;
   RECT 23.18 345.42 157.32 347.13 ;
   RECT 23.18 347.13 157.32 348.84 ;
   RECT 23.18 348.84 157.32 350.55 ;
   RECT 23.18 350.55 157.32 352.26 ;
   RECT 23.18 352.26 157.32 353.97 ;
   RECT 23.18 353.97 157.32 355.68 ;
   RECT 23.18 355.68 157.32 357.39 ;
   RECT 0.0 357.39 157.32 359.1 ;
   RECT 0.0 359.1 157.32 360.81 ;
   RECT 0.0 360.81 157.32 362.52 ;
   RECT 0.0 362.52 157.32 364.23 ;
   RECT 0.0 364.23 157.32 365.94 ;
   RECT 0.0 365.94 157.32 367.65 ;
   RECT 0.0 367.65 157.32 369.36 ;
   RECT 0.0 369.36 157.32 371.07 ;
   RECT 0.0 371.07 157.32 372.78 ;
   RECT 0.0 372.78 157.32 374.49 ;
   RECT 0.0 374.49 157.32 376.2 ;
   RECT 0.0 376.2 157.32 377.91 ;
   RECT 0.0 377.91 157.32 379.62 ;
   RECT 0.0 379.62 157.32 381.33 ;
   RECT 0.0 381.33 157.32 383.04 ;
   RECT 0.0 383.04 157.32 384.75 ;
   RECT 0.0 384.75 157.32 386.46 ;
   RECT 23.18 386.46 157.32 388.17 ;
   RECT 23.18 388.17 157.32 389.88 ;
   RECT 23.18 389.88 157.32 391.59 ;
   RECT 23.18 391.59 157.32 393.3 ;
   RECT 23.18 393.3 157.32 395.01 ;
   RECT 23.18 395.01 157.32 396.72 ;
   RECT 23.18 396.72 157.32 398.43 ;
   RECT 23.18 398.43 157.32 400.14 ;
   RECT 23.18 400.14 157.32 401.85 ;
   RECT 23.18 401.85 157.32 403.56 ;
   RECT 23.18 403.56 157.32 405.27 ;
   RECT 23.18 405.27 157.32 406.98 ;
   RECT 23.18 406.98 157.32 408.69 ;
   RECT 23.18 408.69 157.32 410.4 ;
   RECT 23.18 410.4 157.32 412.11 ;
   RECT 23.18 412.11 157.32 413.82 ;
   RECT 23.18 413.82 157.32 415.53 ;
   RECT 23.18 415.53 157.32 417.24 ;
   RECT 23.18 417.24 157.32 418.95 ;
   RECT 23.18 418.95 157.32 420.66 ;
   RECT 23.18 420.66 157.32 422.37 ;
   RECT 23.18 422.37 157.32 424.08 ;
   RECT 23.18 424.08 157.32 425.79 ;
   RECT 23.18 425.79 157.32 427.5 ;
   RECT 23.18 427.5 157.32 429.21 ;
   RECT 23.18 429.21 157.32 430.92 ;
   RECT 23.18 430.92 157.32 432.63 ;
   RECT 23.18 432.63 157.32 434.34 ;
   RECT 23.18 434.34 157.32 436.05 ;
   RECT 23.18 436.05 157.32 437.76 ;
   RECT 23.18 437.76 157.32 439.47 ;
   RECT 23.18 439.47 157.32 441.18 ;
   RECT 23.18 441.18 157.32 442.89 ;
   RECT 23.18 442.89 157.32 444.6 ;
   RECT 23.18 444.6 157.32 446.31 ;
   RECT 23.18 446.31 157.32 448.02 ;
   RECT 23.18 448.02 157.32 449.73 ;
   RECT 23.18 449.73 157.32 451.44 ;
   RECT 23.18 451.44 157.32 453.15 ;
   RECT 23.18 453.15 157.32 454.86 ;
   RECT 23.18 454.86 157.32 456.57 ;
   RECT 23.18 456.57 157.32 458.28 ;
   RECT 23.18 458.28 157.32 459.99 ;
   RECT 23.18 459.99 157.32 461.7 ;
   RECT 23.18 461.7 157.32 463.41 ;
   RECT 23.18 463.41 157.32 465.12 ;
   RECT 23.18 465.12 157.32 466.83 ;
   RECT 23.18 466.83 157.32 468.54 ;
   RECT 23.18 468.54 157.32 470.25 ;
   RECT 23.18 470.25 157.32 471.96 ;
   RECT 23.18 471.96 157.32 473.67 ;
   RECT 23.18 473.67 157.32 475.38 ;
   RECT 23.18 475.38 157.32 477.09 ;
   RECT 23.18 477.09 157.32 478.8 ;
   RECT 23.18 478.8 157.32 480.51 ;
   RECT 23.18 480.51 157.32 482.22 ;
   RECT 23.18 482.22 157.32 483.93 ;
   RECT 23.18 483.93 157.32 485.64 ;
   RECT 23.18 485.64 157.32 487.35 ;
   RECT 23.18 487.35 157.32 489.06 ;
   RECT 23.18 489.06 157.32 490.77 ;
   RECT 23.18 490.77 157.32 492.48 ;
   RECT 23.18 492.48 157.32 494.19 ;
   RECT 23.18 494.19 157.32 495.9 ;
   RECT 23.18 495.9 157.32 497.61 ;
   RECT 23.18 497.61 157.32 499.32 ;
   RECT 23.18 499.32 157.32 501.03 ;
   RECT 23.18 501.03 157.32 502.74 ;
   RECT 23.18 502.74 157.32 504.45 ;
   RECT 23.18 504.45 157.32 506.16 ;
   RECT 23.18 506.16 157.32 507.87 ;
   RECT 23.18 507.87 157.32 509.58 ;
   RECT 23.18 509.58 157.32 511.29 ;
   RECT 23.18 511.29 157.32 513.0 ;
   RECT 23.18 513.0 157.32 514.71 ;
   RECT 23.18 514.71 157.32 516.42 ;
   RECT 23.18 516.42 157.32 518.13 ;
   RECT 23.18 518.13 157.32 519.84 ;
   RECT 23.18 519.84 157.32 521.55 ;
   RECT 23.18 521.55 157.32 523.26 ;
   RECT 23.18 523.26 157.32 524.97 ;
   RECT 23.18 524.97 157.32 526.68 ;
   RECT 23.18 526.68 157.32 528.39 ;
   RECT 23.18 528.39 157.32 530.1 ;
   RECT 23.18 530.1 157.32 531.81 ;
   RECT 23.18 531.81 157.32 533.52 ;
   RECT 23.18 533.52 157.32 535.23 ;
   RECT 23.18 535.23 157.32 536.94 ;
   RECT 23.18 536.94 157.32 538.65 ;
   RECT 23.18 538.65 157.32 540.36 ;
   RECT 23.18 540.36 157.32 542.07 ;
   RECT 23.18 542.07 157.32 543.78 ;
   RECT 23.18 543.78 157.32 545.49 ;
   RECT 23.18 545.49 157.32 547.2 ;
   RECT 23.18 547.2 157.32 548.91 ;
   RECT 23.18 548.91 157.32 550.62 ;
   RECT 23.18 550.62 157.32 552.33 ;
   RECT 23.18 552.33 157.32 554.04 ;
   RECT 23.18 554.04 157.32 555.75 ;
   RECT 23.18 555.75 157.32 557.46 ;
   RECT 23.18 557.46 157.32 559.17 ;
   RECT 23.18 559.17 157.32 560.88 ;
   RECT 23.18 560.88 157.32 562.59 ;
   RECT 23.18 562.59 157.32 564.3 ;
   RECT 23.18 564.3 157.32 566.01 ;
   RECT 23.18 566.01 157.32 567.72 ;
   RECT 23.18 567.72 157.32 569.43 ;
   RECT 23.18 569.43 157.32 571.14 ;
   RECT 23.18 571.14 157.32 572.85 ;
   RECT 23.18 572.85 157.32 574.56 ;
   RECT 23.18 574.56 157.32 576.27 ;
   RECT 23.18 576.27 157.32 577.98 ;
   RECT 23.18 577.98 157.32 579.69 ;
   RECT 23.18 579.69 157.32 581.4 ;
   RECT 23.18 581.4 157.32 583.11 ;
   RECT 23.18 583.11 157.32 584.82 ;
   RECT 23.18 584.82 157.32 586.53 ;
   RECT 23.18 586.53 157.32 588.24 ;
   RECT 23.18 588.24 157.32 589.95 ;
   RECT 23.18 589.95 157.32 591.66 ;
   RECT 23.18 591.66 157.32 593.37 ;
   RECT 23.18 593.37 157.32 595.08 ;
   RECT 23.18 595.08 157.32 596.79 ;
   RECT 23.18 596.79 157.32 598.5 ;
   RECT 23.18 598.5 157.32 600.21 ;
   RECT 23.18 600.21 157.32 601.92 ;
   RECT 23.18 601.92 157.32 603.63 ;
   RECT 23.18 603.63 157.32 605.34 ;
   RECT 23.18 605.34 157.32 607.05 ;
   RECT 23.18 607.05 157.32 608.76 ;
   RECT 23.18 608.76 157.32 610.47 ;
   RECT 23.18 610.47 157.32 612.18 ;
   RECT 23.18 612.18 157.32 613.89 ;
   RECT 23.18 613.89 157.32 615.6 ;
   RECT 23.18 615.6 157.32 617.31 ;
   RECT 23.18 617.31 157.32 619.02 ;
   RECT 23.18 619.02 157.32 620.73 ;
   RECT 23.18 620.73 157.32 622.44 ;
   RECT 23.18 622.44 157.32 624.15 ;
   RECT 23.18 624.15 157.32 625.86 ;
   RECT 23.18 625.86 157.32 627.57 ;
   RECT 23.18 627.57 157.32 629.28 ;
   RECT 23.18 629.28 157.32 630.99 ;
   RECT 23.18 630.99 157.32 632.7 ;
   RECT 23.18 632.7 157.32 634.41 ;
   RECT 23.18 634.41 157.32 636.12 ;
   RECT 23.18 636.12 157.32 637.83 ;
   RECT 23.18 637.83 157.32 639.54 ;
   RECT 23.18 639.54 157.32 641.25 ;
   RECT 23.18 641.25 157.32 642.96 ;
   RECT 23.18 642.96 157.32 644.67 ;
   RECT 23.18 644.67 157.32 646.38 ;
   RECT 23.18 646.38 157.32 648.09 ;
   RECT 23.18 648.09 157.32 649.8 ;
   RECT 23.18 649.8 157.32 651.51 ;
   RECT 23.18 651.51 157.32 653.22 ;
   RECT 23.18 653.22 157.32 654.93 ;
   RECT 23.18 654.93 157.32 656.64 ;
   RECT 23.18 656.64 157.32 658.35 ;
   RECT 23.18 658.35 157.32 660.06 ;
   RECT 23.18 660.06 157.32 661.77 ;
   RECT 23.18 661.77 157.32 663.48 ;
   RECT 23.18 663.48 157.32 665.19 ;
   RECT 23.18 665.19 157.32 666.9 ;
   RECT 23.18 666.9 157.32 668.61 ;
   RECT 23.18 668.61 157.32 670.32 ;
   RECT 23.18 670.32 157.32 672.03 ;
   RECT 23.18 672.03 157.32 673.74 ;
   RECT 23.18 673.74 157.32 675.45 ;
   RECT 23.18 675.45 157.32 677.16 ;
   RECT 23.18 677.16 157.32 678.87 ;
   RECT 23.18 678.87 157.32 680.58 ;
   RECT 23.18 680.58 157.32 682.29 ;
   RECT 23.18 682.29 157.32 684.0 ;
   RECT 23.18 684.0 157.32 685.71 ;
   RECT 23.18 685.71 157.32 687.42 ;
   RECT 23.18 687.42 157.32 689.13 ;
   RECT 23.18 689.13 157.32 690.84 ;
   RECT 23.18 690.84 157.32 692.55 ;
   RECT 23.18 692.55 157.32 694.26 ;
   RECT 23.18 694.26 157.32 695.97 ;
   RECT 23.18 695.97 157.32 697.68 ;
   RECT 23.18 697.68 157.32 699.39 ;
   RECT 23.18 699.39 157.32 701.1 ;
   RECT 23.18 701.1 157.32 702.81 ;
   RECT 23.18 702.81 157.32 704.52 ;
   RECT 23.18 704.52 157.32 706.23 ;
   RECT 23.18 706.23 157.32 707.94 ;
   RECT 23.18 707.94 157.32 709.65 ;
   RECT 23.18 709.65 157.32 711.36 ;
   RECT 23.18 711.36 157.32 713.07 ;
   RECT 23.18 713.07 157.32 714.78 ;
   RECT 23.18 714.78 157.32 716.49 ;
   RECT 23.18 716.49 157.32 718.2 ;
   RECT 23.18 718.2 157.32 719.91 ;
   RECT 23.18 719.91 157.32 721.62 ;
   RECT 23.18 721.62 157.32 723.33 ;
   RECT 23.18 723.33 157.32 725.04 ;
   RECT 23.18 725.04 157.32 726.75 ;
   RECT 23.18 726.75 157.32 728.46 ;
   RECT 23.18 728.46 157.32 730.17 ;
   RECT 23.18 730.17 157.32 731.88 ;
   RECT 23.18 731.88 157.32 733.59 ;
   RECT 23.18 733.59 157.32 735.3 ;
   RECT 23.18 735.3 157.32 737.01 ;
   RECT 23.18 737.01 157.32 738.72 ;
   RECT 23.18 738.72 157.32 740.43 ;
   RECT 23.18 740.43 157.32 742.14 ;
   RECT 23.18 742.14 157.32 743.85 ;
   RECT 23.18 743.85 157.32 745.56 ;
   RECT 23.18 745.56 157.32 747.27 ;
   RECT 23.18 747.27 157.32 748.98 ;
   RECT 23.18 748.98 157.32 750.69 ;
   RECT 23.18 750.69 157.32 752.4 ;
   RECT 23.18 752.4 157.32 754.11 ;
   RECT 23.18 754.11 157.32 755.82 ;
  LAYER via2 ;
   RECT 23.18 0.0 157.32 1.71 ;
   RECT 23.18 1.71 157.32 3.42 ;
   RECT 23.18 3.42 157.32 5.13 ;
   RECT 23.18 5.13 157.32 6.84 ;
   RECT 23.18 6.84 157.32 8.55 ;
   RECT 23.18 8.55 157.32 10.26 ;
   RECT 23.18 10.26 157.32 11.97 ;
   RECT 23.18 11.97 157.32 13.68 ;
   RECT 23.18 13.68 157.32 15.39 ;
   RECT 23.18 15.39 157.32 17.1 ;
   RECT 23.18 17.1 157.32 18.81 ;
   RECT 23.18 18.81 157.32 20.52 ;
   RECT 23.18 20.52 157.32 22.23 ;
   RECT 23.18 22.23 157.32 23.94 ;
   RECT 23.18 23.94 157.32 25.65 ;
   RECT 23.18 25.65 157.32 27.36 ;
   RECT 23.18 27.36 157.32 29.07 ;
   RECT 23.18 29.07 157.32 30.78 ;
   RECT 23.18 30.78 157.32 32.49 ;
   RECT 23.18 32.49 157.32 34.2 ;
   RECT 23.18 34.2 157.32 35.91 ;
   RECT 23.18 35.91 157.32 37.62 ;
   RECT 23.18 37.62 157.32 39.33 ;
   RECT 23.18 39.33 157.32 41.04 ;
   RECT 23.18 41.04 157.32 42.75 ;
   RECT 23.18 42.75 157.32 44.46 ;
   RECT 23.18 44.46 157.32 46.17 ;
   RECT 23.18 46.17 157.32 47.88 ;
   RECT 23.18 47.88 157.32 49.59 ;
   RECT 23.18 49.59 157.32 51.3 ;
   RECT 23.18 51.3 157.32 53.01 ;
   RECT 23.18 53.01 157.32 54.72 ;
   RECT 23.18 54.72 157.32 56.43 ;
   RECT 23.18 56.43 157.32 58.14 ;
   RECT 23.18 58.14 157.32 59.85 ;
   RECT 23.18 59.85 157.32 61.56 ;
   RECT 23.18 61.56 157.32 63.27 ;
   RECT 23.18 63.27 157.32 64.98 ;
   RECT 23.18 64.98 157.32 66.69 ;
   RECT 23.18 66.69 157.32 68.4 ;
   RECT 23.18 68.4 157.32 70.11 ;
   RECT 23.18 70.11 157.32 71.82 ;
   RECT 23.18 71.82 157.32 73.53 ;
   RECT 23.18 73.53 157.32 75.24 ;
   RECT 23.18 75.24 157.32 76.95 ;
   RECT 23.18 76.95 157.32 78.66 ;
   RECT 23.18 78.66 157.32 80.37 ;
   RECT 23.18 80.37 157.32 82.08 ;
   RECT 23.18 82.08 157.32 83.79 ;
   RECT 23.18 83.79 157.32 85.5 ;
   RECT 23.18 85.5 157.32 87.21 ;
   RECT 23.18 87.21 157.32 88.92 ;
   RECT 23.18 88.92 157.32 90.63 ;
   RECT 23.18 90.63 157.32 92.34 ;
   RECT 23.18 92.34 157.32 94.05 ;
   RECT 23.18 94.05 157.32 95.76 ;
   RECT 23.18 95.76 157.32 97.47 ;
   RECT 23.18 97.47 157.32 99.18 ;
   RECT 23.18 99.18 157.32 100.89 ;
   RECT 23.18 100.89 157.32 102.6 ;
   RECT 23.18 102.6 157.32 104.31 ;
   RECT 23.18 104.31 157.32 106.02 ;
   RECT 23.18 106.02 157.32 107.73 ;
   RECT 23.18 107.73 157.32 109.44 ;
   RECT 23.18 109.44 157.32 111.15 ;
   RECT 23.18 111.15 157.32 112.86 ;
   RECT 23.18 112.86 157.32 114.57 ;
   RECT 23.18 114.57 157.32 116.28 ;
   RECT 23.18 116.28 157.32 117.99 ;
   RECT 23.18 117.99 157.32 119.7 ;
   RECT 23.18 119.7 157.32 121.41 ;
   RECT 23.18 121.41 157.32 123.12 ;
   RECT 23.18 123.12 157.32 124.83 ;
   RECT 23.18 124.83 157.32 126.54 ;
   RECT 23.18 126.54 157.32 128.25 ;
   RECT 23.18 128.25 157.32 129.96 ;
   RECT 23.18 129.96 157.32 131.67 ;
   RECT 23.18 131.67 157.32 133.38 ;
   RECT 23.18 133.38 157.32 135.09 ;
   RECT 23.18 135.09 157.32 136.8 ;
   RECT 23.18 136.8 157.32 138.51 ;
   RECT 23.18 138.51 157.32 140.22 ;
   RECT 23.18 140.22 157.32 141.93 ;
   RECT 23.18 141.93 157.32 143.64 ;
   RECT 23.18 143.64 157.32 145.35 ;
   RECT 23.18 145.35 157.32 147.06 ;
   RECT 23.18 147.06 157.32 148.77 ;
   RECT 23.18 148.77 157.32 150.48 ;
   RECT 23.18 150.48 157.32 152.19 ;
   RECT 23.18 152.19 157.32 153.9 ;
   RECT 23.18 153.9 157.32 155.61 ;
   RECT 23.18 155.61 157.32 157.32 ;
   RECT 23.18 157.32 157.32 159.03 ;
   RECT 23.18 159.03 157.32 160.74 ;
   RECT 23.18 160.74 157.32 162.45 ;
   RECT 23.18 162.45 157.32 164.16 ;
   RECT 23.18 164.16 157.32 165.87 ;
   RECT 23.18 165.87 157.32 167.58 ;
   RECT 23.18 167.58 157.32 169.29 ;
   RECT 23.18 169.29 157.32 171.0 ;
   RECT 23.18 171.0 157.32 172.71 ;
   RECT 23.18 172.71 157.32 174.42 ;
   RECT 23.18 174.42 157.32 176.13 ;
   RECT 23.18 176.13 157.32 177.84 ;
   RECT 23.18 177.84 157.32 179.55 ;
   RECT 23.18 179.55 157.32 181.26 ;
   RECT 23.18 181.26 157.32 182.97 ;
   RECT 23.18 182.97 157.32 184.68 ;
   RECT 23.18 184.68 157.32 186.39 ;
   RECT 23.18 186.39 157.32 188.1 ;
   RECT 23.18 188.1 157.32 189.81 ;
   RECT 23.18 189.81 157.32 191.52 ;
   RECT 23.18 191.52 157.32 193.23 ;
   RECT 23.18 193.23 157.32 194.94 ;
   RECT 23.18 194.94 157.32 196.65 ;
   RECT 23.18 196.65 157.32 198.36 ;
   RECT 23.18 198.36 157.32 200.07 ;
   RECT 23.18 200.07 157.32 201.78 ;
   RECT 23.18 201.78 157.32 203.49 ;
   RECT 23.18 203.49 157.32 205.2 ;
   RECT 23.18 205.2 157.32 206.91 ;
   RECT 23.18 206.91 157.32 208.62 ;
   RECT 23.18 208.62 157.32 210.33 ;
   RECT 23.18 210.33 157.32 212.04 ;
   RECT 23.18 212.04 157.32 213.75 ;
   RECT 23.18 213.75 157.32 215.46 ;
   RECT 23.18 215.46 157.32 217.17 ;
   RECT 23.18 217.17 157.32 218.88 ;
   RECT 23.18 218.88 157.32 220.59 ;
   RECT 23.18 220.59 157.32 222.3 ;
   RECT 23.18 222.3 157.32 224.01 ;
   RECT 23.18 224.01 157.32 225.72 ;
   RECT 23.18 225.72 157.32 227.43 ;
   RECT 23.18 227.43 157.32 229.14 ;
   RECT 23.18 229.14 157.32 230.85 ;
   RECT 23.18 230.85 157.32 232.56 ;
   RECT 23.18 232.56 157.32 234.27 ;
   RECT 23.18 234.27 157.32 235.98 ;
   RECT 23.18 235.98 157.32 237.69 ;
   RECT 23.18 237.69 157.32 239.4 ;
   RECT 23.18 239.4 157.32 241.11 ;
   RECT 23.18 241.11 157.32 242.82 ;
   RECT 23.18 242.82 157.32 244.53 ;
   RECT 23.18 244.53 157.32 246.24 ;
   RECT 23.18 246.24 157.32 247.95 ;
   RECT 23.18 247.95 157.32 249.66 ;
   RECT 23.18 249.66 157.32 251.37 ;
   RECT 23.18 251.37 157.32 253.08 ;
   RECT 23.18 253.08 157.32 254.79 ;
   RECT 23.18 254.79 157.32 256.5 ;
   RECT 23.18 256.5 157.32 258.21 ;
   RECT 23.18 258.21 157.32 259.92 ;
   RECT 23.18 259.92 157.32 261.63 ;
   RECT 23.18 261.63 157.32 263.34 ;
   RECT 23.18 263.34 157.32 265.05 ;
   RECT 23.18 265.05 157.32 266.76 ;
   RECT 23.18 266.76 157.32 268.47 ;
   RECT 23.18 268.47 157.32 270.18 ;
   RECT 23.18 270.18 157.32 271.89 ;
   RECT 23.18 271.89 157.32 273.6 ;
   RECT 23.18 273.6 157.32 275.31 ;
   RECT 23.18 275.31 157.32 277.02 ;
   RECT 23.18 277.02 157.32 278.73 ;
   RECT 23.18 278.73 157.32 280.44 ;
   RECT 23.18 280.44 157.32 282.15 ;
   RECT 23.18 282.15 157.32 283.86 ;
   RECT 23.18 283.86 157.32 285.57 ;
   RECT 23.18 285.57 157.32 287.28 ;
   RECT 23.18 287.28 157.32 288.99 ;
   RECT 23.18 288.99 157.32 290.7 ;
   RECT 23.18 290.7 157.32 292.41 ;
   RECT 23.18 292.41 157.32 294.12 ;
   RECT 23.18 294.12 157.32 295.83 ;
   RECT 23.18 295.83 157.32 297.54 ;
   RECT 23.18 297.54 157.32 299.25 ;
   RECT 23.18 299.25 157.32 300.96 ;
   RECT 23.18 300.96 157.32 302.67 ;
   RECT 23.18 302.67 157.32 304.38 ;
   RECT 23.18 304.38 157.32 306.09 ;
   RECT 23.18 306.09 157.32 307.8 ;
   RECT 23.18 307.8 157.32 309.51 ;
   RECT 23.18 309.51 157.32 311.22 ;
   RECT 23.18 311.22 157.32 312.93 ;
   RECT 23.18 312.93 157.32 314.64 ;
   RECT 23.18 314.64 157.32 316.35 ;
   RECT 23.18 316.35 157.32 318.06 ;
   RECT 23.18 318.06 157.32 319.77 ;
   RECT 23.18 319.77 157.32 321.48 ;
   RECT 23.18 321.48 157.32 323.19 ;
   RECT 23.18 323.19 157.32 324.9 ;
   RECT 23.18 324.9 157.32 326.61 ;
   RECT 23.18 326.61 157.32 328.32 ;
   RECT 23.18 328.32 157.32 330.03 ;
   RECT 23.18 330.03 157.32 331.74 ;
   RECT 23.18 331.74 157.32 333.45 ;
   RECT 23.18 333.45 157.32 335.16 ;
   RECT 23.18 335.16 157.32 336.87 ;
   RECT 23.18 336.87 157.32 338.58 ;
   RECT 23.18 338.58 157.32 340.29 ;
   RECT 23.18 340.29 157.32 342.0 ;
   RECT 23.18 342.0 157.32 343.71 ;
   RECT 23.18 343.71 157.32 345.42 ;
   RECT 23.18 345.42 157.32 347.13 ;
   RECT 23.18 347.13 157.32 348.84 ;
   RECT 23.18 348.84 157.32 350.55 ;
   RECT 23.18 350.55 157.32 352.26 ;
   RECT 23.18 352.26 157.32 353.97 ;
   RECT 23.18 353.97 157.32 355.68 ;
   RECT 23.18 355.68 157.32 357.39 ;
   RECT 0.0 357.39 157.32 359.1 ;
   RECT 0.0 359.1 157.32 360.81 ;
   RECT 0.0 360.81 157.32 362.52 ;
   RECT 0.0 362.52 157.32 364.23 ;
   RECT 0.0 364.23 157.32 365.94 ;
   RECT 0.0 365.94 157.32 367.65 ;
   RECT 0.0 367.65 157.32 369.36 ;
   RECT 0.0 369.36 157.32 371.07 ;
   RECT 0.0 371.07 157.32 372.78 ;
   RECT 0.0 372.78 157.32 374.49 ;
   RECT 0.0 374.49 157.32 376.2 ;
   RECT 0.0 376.2 157.32 377.91 ;
   RECT 0.0 377.91 157.32 379.62 ;
   RECT 0.0 379.62 157.32 381.33 ;
   RECT 0.0 381.33 157.32 383.04 ;
   RECT 0.0 383.04 157.32 384.75 ;
   RECT 0.0 384.75 157.32 386.46 ;
   RECT 23.18 386.46 157.32 388.17 ;
   RECT 23.18 388.17 157.32 389.88 ;
   RECT 23.18 389.88 157.32 391.59 ;
   RECT 23.18 391.59 157.32 393.3 ;
   RECT 23.18 393.3 157.32 395.01 ;
   RECT 23.18 395.01 157.32 396.72 ;
   RECT 23.18 396.72 157.32 398.43 ;
   RECT 23.18 398.43 157.32 400.14 ;
   RECT 23.18 400.14 157.32 401.85 ;
   RECT 23.18 401.85 157.32 403.56 ;
   RECT 23.18 403.56 157.32 405.27 ;
   RECT 23.18 405.27 157.32 406.98 ;
   RECT 23.18 406.98 157.32 408.69 ;
   RECT 23.18 408.69 157.32 410.4 ;
   RECT 23.18 410.4 157.32 412.11 ;
   RECT 23.18 412.11 157.32 413.82 ;
   RECT 23.18 413.82 157.32 415.53 ;
   RECT 23.18 415.53 157.32 417.24 ;
   RECT 23.18 417.24 157.32 418.95 ;
   RECT 23.18 418.95 157.32 420.66 ;
   RECT 23.18 420.66 157.32 422.37 ;
   RECT 23.18 422.37 157.32 424.08 ;
   RECT 23.18 424.08 157.32 425.79 ;
   RECT 23.18 425.79 157.32 427.5 ;
   RECT 23.18 427.5 157.32 429.21 ;
   RECT 23.18 429.21 157.32 430.92 ;
   RECT 23.18 430.92 157.32 432.63 ;
   RECT 23.18 432.63 157.32 434.34 ;
   RECT 23.18 434.34 157.32 436.05 ;
   RECT 23.18 436.05 157.32 437.76 ;
   RECT 23.18 437.76 157.32 439.47 ;
   RECT 23.18 439.47 157.32 441.18 ;
   RECT 23.18 441.18 157.32 442.89 ;
   RECT 23.18 442.89 157.32 444.6 ;
   RECT 23.18 444.6 157.32 446.31 ;
   RECT 23.18 446.31 157.32 448.02 ;
   RECT 23.18 448.02 157.32 449.73 ;
   RECT 23.18 449.73 157.32 451.44 ;
   RECT 23.18 451.44 157.32 453.15 ;
   RECT 23.18 453.15 157.32 454.86 ;
   RECT 23.18 454.86 157.32 456.57 ;
   RECT 23.18 456.57 157.32 458.28 ;
   RECT 23.18 458.28 157.32 459.99 ;
   RECT 23.18 459.99 157.32 461.7 ;
   RECT 23.18 461.7 157.32 463.41 ;
   RECT 23.18 463.41 157.32 465.12 ;
   RECT 23.18 465.12 157.32 466.83 ;
   RECT 23.18 466.83 157.32 468.54 ;
   RECT 23.18 468.54 157.32 470.25 ;
   RECT 23.18 470.25 157.32 471.96 ;
   RECT 23.18 471.96 157.32 473.67 ;
   RECT 23.18 473.67 157.32 475.38 ;
   RECT 23.18 475.38 157.32 477.09 ;
   RECT 23.18 477.09 157.32 478.8 ;
   RECT 23.18 478.8 157.32 480.51 ;
   RECT 23.18 480.51 157.32 482.22 ;
   RECT 23.18 482.22 157.32 483.93 ;
   RECT 23.18 483.93 157.32 485.64 ;
   RECT 23.18 485.64 157.32 487.35 ;
   RECT 23.18 487.35 157.32 489.06 ;
   RECT 23.18 489.06 157.32 490.77 ;
   RECT 23.18 490.77 157.32 492.48 ;
   RECT 23.18 492.48 157.32 494.19 ;
   RECT 23.18 494.19 157.32 495.9 ;
   RECT 23.18 495.9 157.32 497.61 ;
   RECT 23.18 497.61 157.32 499.32 ;
   RECT 23.18 499.32 157.32 501.03 ;
   RECT 23.18 501.03 157.32 502.74 ;
   RECT 23.18 502.74 157.32 504.45 ;
   RECT 23.18 504.45 157.32 506.16 ;
   RECT 23.18 506.16 157.32 507.87 ;
   RECT 23.18 507.87 157.32 509.58 ;
   RECT 23.18 509.58 157.32 511.29 ;
   RECT 23.18 511.29 157.32 513.0 ;
   RECT 23.18 513.0 157.32 514.71 ;
   RECT 23.18 514.71 157.32 516.42 ;
   RECT 23.18 516.42 157.32 518.13 ;
   RECT 23.18 518.13 157.32 519.84 ;
   RECT 23.18 519.84 157.32 521.55 ;
   RECT 23.18 521.55 157.32 523.26 ;
   RECT 23.18 523.26 157.32 524.97 ;
   RECT 23.18 524.97 157.32 526.68 ;
   RECT 23.18 526.68 157.32 528.39 ;
   RECT 23.18 528.39 157.32 530.1 ;
   RECT 23.18 530.1 157.32 531.81 ;
   RECT 23.18 531.81 157.32 533.52 ;
   RECT 23.18 533.52 157.32 535.23 ;
   RECT 23.18 535.23 157.32 536.94 ;
   RECT 23.18 536.94 157.32 538.65 ;
   RECT 23.18 538.65 157.32 540.36 ;
   RECT 23.18 540.36 157.32 542.07 ;
   RECT 23.18 542.07 157.32 543.78 ;
   RECT 23.18 543.78 157.32 545.49 ;
   RECT 23.18 545.49 157.32 547.2 ;
   RECT 23.18 547.2 157.32 548.91 ;
   RECT 23.18 548.91 157.32 550.62 ;
   RECT 23.18 550.62 157.32 552.33 ;
   RECT 23.18 552.33 157.32 554.04 ;
   RECT 23.18 554.04 157.32 555.75 ;
   RECT 23.18 555.75 157.32 557.46 ;
   RECT 23.18 557.46 157.32 559.17 ;
   RECT 23.18 559.17 157.32 560.88 ;
   RECT 23.18 560.88 157.32 562.59 ;
   RECT 23.18 562.59 157.32 564.3 ;
   RECT 23.18 564.3 157.32 566.01 ;
   RECT 23.18 566.01 157.32 567.72 ;
   RECT 23.18 567.72 157.32 569.43 ;
   RECT 23.18 569.43 157.32 571.14 ;
   RECT 23.18 571.14 157.32 572.85 ;
   RECT 23.18 572.85 157.32 574.56 ;
   RECT 23.18 574.56 157.32 576.27 ;
   RECT 23.18 576.27 157.32 577.98 ;
   RECT 23.18 577.98 157.32 579.69 ;
   RECT 23.18 579.69 157.32 581.4 ;
   RECT 23.18 581.4 157.32 583.11 ;
   RECT 23.18 583.11 157.32 584.82 ;
   RECT 23.18 584.82 157.32 586.53 ;
   RECT 23.18 586.53 157.32 588.24 ;
   RECT 23.18 588.24 157.32 589.95 ;
   RECT 23.18 589.95 157.32 591.66 ;
   RECT 23.18 591.66 157.32 593.37 ;
   RECT 23.18 593.37 157.32 595.08 ;
   RECT 23.18 595.08 157.32 596.79 ;
   RECT 23.18 596.79 157.32 598.5 ;
   RECT 23.18 598.5 157.32 600.21 ;
   RECT 23.18 600.21 157.32 601.92 ;
   RECT 23.18 601.92 157.32 603.63 ;
   RECT 23.18 603.63 157.32 605.34 ;
   RECT 23.18 605.34 157.32 607.05 ;
   RECT 23.18 607.05 157.32 608.76 ;
   RECT 23.18 608.76 157.32 610.47 ;
   RECT 23.18 610.47 157.32 612.18 ;
   RECT 23.18 612.18 157.32 613.89 ;
   RECT 23.18 613.89 157.32 615.6 ;
   RECT 23.18 615.6 157.32 617.31 ;
   RECT 23.18 617.31 157.32 619.02 ;
   RECT 23.18 619.02 157.32 620.73 ;
   RECT 23.18 620.73 157.32 622.44 ;
   RECT 23.18 622.44 157.32 624.15 ;
   RECT 23.18 624.15 157.32 625.86 ;
   RECT 23.18 625.86 157.32 627.57 ;
   RECT 23.18 627.57 157.32 629.28 ;
   RECT 23.18 629.28 157.32 630.99 ;
   RECT 23.18 630.99 157.32 632.7 ;
   RECT 23.18 632.7 157.32 634.41 ;
   RECT 23.18 634.41 157.32 636.12 ;
   RECT 23.18 636.12 157.32 637.83 ;
   RECT 23.18 637.83 157.32 639.54 ;
   RECT 23.18 639.54 157.32 641.25 ;
   RECT 23.18 641.25 157.32 642.96 ;
   RECT 23.18 642.96 157.32 644.67 ;
   RECT 23.18 644.67 157.32 646.38 ;
   RECT 23.18 646.38 157.32 648.09 ;
   RECT 23.18 648.09 157.32 649.8 ;
   RECT 23.18 649.8 157.32 651.51 ;
   RECT 23.18 651.51 157.32 653.22 ;
   RECT 23.18 653.22 157.32 654.93 ;
   RECT 23.18 654.93 157.32 656.64 ;
   RECT 23.18 656.64 157.32 658.35 ;
   RECT 23.18 658.35 157.32 660.06 ;
   RECT 23.18 660.06 157.32 661.77 ;
   RECT 23.18 661.77 157.32 663.48 ;
   RECT 23.18 663.48 157.32 665.19 ;
   RECT 23.18 665.19 157.32 666.9 ;
   RECT 23.18 666.9 157.32 668.61 ;
   RECT 23.18 668.61 157.32 670.32 ;
   RECT 23.18 670.32 157.32 672.03 ;
   RECT 23.18 672.03 157.32 673.74 ;
   RECT 23.18 673.74 157.32 675.45 ;
   RECT 23.18 675.45 157.32 677.16 ;
   RECT 23.18 677.16 157.32 678.87 ;
   RECT 23.18 678.87 157.32 680.58 ;
   RECT 23.18 680.58 157.32 682.29 ;
   RECT 23.18 682.29 157.32 684.0 ;
   RECT 23.18 684.0 157.32 685.71 ;
   RECT 23.18 685.71 157.32 687.42 ;
   RECT 23.18 687.42 157.32 689.13 ;
   RECT 23.18 689.13 157.32 690.84 ;
   RECT 23.18 690.84 157.32 692.55 ;
   RECT 23.18 692.55 157.32 694.26 ;
   RECT 23.18 694.26 157.32 695.97 ;
   RECT 23.18 695.97 157.32 697.68 ;
   RECT 23.18 697.68 157.32 699.39 ;
   RECT 23.18 699.39 157.32 701.1 ;
   RECT 23.18 701.1 157.32 702.81 ;
   RECT 23.18 702.81 157.32 704.52 ;
   RECT 23.18 704.52 157.32 706.23 ;
   RECT 23.18 706.23 157.32 707.94 ;
   RECT 23.18 707.94 157.32 709.65 ;
   RECT 23.18 709.65 157.32 711.36 ;
   RECT 23.18 711.36 157.32 713.07 ;
   RECT 23.18 713.07 157.32 714.78 ;
   RECT 23.18 714.78 157.32 716.49 ;
   RECT 23.18 716.49 157.32 718.2 ;
   RECT 23.18 718.2 157.32 719.91 ;
   RECT 23.18 719.91 157.32 721.62 ;
   RECT 23.18 721.62 157.32 723.33 ;
   RECT 23.18 723.33 157.32 725.04 ;
   RECT 23.18 725.04 157.32 726.75 ;
   RECT 23.18 726.75 157.32 728.46 ;
   RECT 23.18 728.46 157.32 730.17 ;
   RECT 23.18 730.17 157.32 731.88 ;
   RECT 23.18 731.88 157.32 733.59 ;
   RECT 23.18 733.59 157.32 735.3 ;
   RECT 23.18 735.3 157.32 737.01 ;
   RECT 23.18 737.01 157.32 738.72 ;
   RECT 23.18 738.72 157.32 740.43 ;
   RECT 23.18 740.43 157.32 742.14 ;
   RECT 23.18 742.14 157.32 743.85 ;
   RECT 23.18 743.85 157.32 745.56 ;
   RECT 23.18 745.56 157.32 747.27 ;
   RECT 23.18 747.27 157.32 748.98 ;
   RECT 23.18 748.98 157.32 750.69 ;
   RECT 23.18 750.69 157.32 752.4 ;
   RECT 23.18 752.4 157.32 754.11 ;
   RECT 23.18 754.11 157.32 755.82 ;
  LAYER metal3 ;
   RECT 23.18 0.0 157.32 1.71 ;
   RECT 23.18 1.71 157.32 3.42 ;
   RECT 23.18 3.42 157.32 5.13 ;
   RECT 23.18 5.13 157.32 6.84 ;
   RECT 23.18 6.84 157.32 8.55 ;
   RECT 23.18 8.55 157.32 10.26 ;
   RECT 23.18 10.26 157.32 11.97 ;
   RECT 23.18 11.97 157.32 13.68 ;
   RECT 23.18 13.68 157.32 15.39 ;
   RECT 23.18 15.39 157.32 17.1 ;
   RECT 23.18 17.1 157.32 18.81 ;
   RECT 23.18 18.81 157.32 20.52 ;
   RECT 23.18 20.52 157.32 22.23 ;
   RECT 23.18 22.23 157.32 23.94 ;
   RECT 23.18 23.94 157.32 25.65 ;
   RECT 23.18 25.65 157.32 27.36 ;
   RECT 23.18 27.36 157.32 29.07 ;
   RECT 23.18 29.07 157.32 30.78 ;
   RECT 23.18 30.78 157.32 32.49 ;
   RECT 23.18 32.49 157.32 34.2 ;
   RECT 23.18 34.2 157.32 35.91 ;
   RECT 23.18 35.91 157.32 37.62 ;
   RECT 23.18 37.62 157.32 39.33 ;
   RECT 23.18 39.33 157.32 41.04 ;
   RECT 23.18 41.04 157.32 42.75 ;
   RECT 23.18 42.75 157.32 44.46 ;
   RECT 23.18 44.46 157.32 46.17 ;
   RECT 23.18 46.17 157.32 47.88 ;
   RECT 23.18 47.88 157.32 49.59 ;
   RECT 23.18 49.59 157.32 51.3 ;
   RECT 23.18 51.3 157.32 53.01 ;
   RECT 23.18 53.01 157.32 54.72 ;
   RECT 23.18 54.72 157.32 56.43 ;
   RECT 23.18 56.43 157.32 58.14 ;
   RECT 23.18 58.14 157.32 59.85 ;
   RECT 23.18 59.85 157.32 61.56 ;
   RECT 23.18 61.56 157.32 63.27 ;
   RECT 23.18 63.27 157.32 64.98 ;
   RECT 23.18 64.98 157.32 66.69 ;
   RECT 23.18 66.69 157.32 68.4 ;
   RECT 23.18 68.4 157.32 70.11 ;
   RECT 23.18 70.11 157.32 71.82 ;
   RECT 23.18 71.82 157.32 73.53 ;
   RECT 23.18 73.53 157.32 75.24 ;
   RECT 23.18 75.24 157.32 76.95 ;
   RECT 23.18 76.95 157.32 78.66 ;
   RECT 23.18 78.66 157.32 80.37 ;
   RECT 23.18 80.37 157.32 82.08 ;
   RECT 23.18 82.08 157.32 83.79 ;
   RECT 23.18 83.79 157.32 85.5 ;
   RECT 23.18 85.5 157.32 87.21 ;
   RECT 23.18 87.21 157.32 88.92 ;
   RECT 23.18 88.92 157.32 90.63 ;
   RECT 23.18 90.63 157.32 92.34 ;
   RECT 23.18 92.34 157.32 94.05 ;
   RECT 23.18 94.05 157.32 95.76 ;
   RECT 23.18 95.76 157.32 97.47 ;
   RECT 23.18 97.47 157.32 99.18 ;
   RECT 23.18 99.18 157.32 100.89 ;
   RECT 23.18 100.89 157.32 102.6 ;
   RECT 23.18 102.6 157.32 104.31 ;
   RECT 23.18 104.31 157.32 106.02 ;
   RECT 23.18 106.02 157.32 107.73 ;
   RECT 23.18 107.73 157.32 109.44 ;
   RECT 23.18 109.44 157.32 111.15 ;
   RECT 23.18 111.15 157.32 112.86 ;
   RECT 23.18 112.86 157.32 114.57 ;
   RECT 23.18 114.57 157.32 116.28 ;
   RECT 23.18 116.28 157.32 117.99 ;
   RECT 23.18 117.99 157.32 119.7 ;
   RECT 23.18 119.7 157.32 121.41 ;
   RECT 23.18 121.41 157.32 123.12 ;
   RECT 23.18 123.12 157.32 124.83 ;
   RECT 23.18 124.83 157.32 126.54 ;
   RECT 23.18 126.54 157.32 128.25 ;
   RECT 23.18 128.25 157.32 129.96 ;
   RECT 23.18 129.96 157.32 131.67 ;
   RECT 23.18 131.67 157.32 133.38 ;
   RECT 23.18 133.38 157.32 135.09 ;
   RECT 23.18 135.09 157.32 136.8 ;
   RECT 23.18 136.8 157.32 138.51 ;
   RECT 23.18 138.51 157.32 140.22 ;
   RECT 23.18 140.22 157.32 141.93 ;
   RECT 23.18 141.93 157.32 143.64 ;
   RECT 23.18 143.64 157.32 145.35 ;
   RECT 23.18 145.35 157.32 147.06 ;
   RECT 23.18 147.06 157.32 148.77 ;
   RECT 23.18 148.77 157.32 150.48 ;
   RECT 23.18 150.48 157.32 152.19 ;
   RECT 23.18 152.19 157.32 153.9 ;
   RECT 23.18 153.9 157.32 155.61 ;
   RECT 23.18 155.61 157.32 157.32 ;
   RECT 23.18 157.32 157.32 159.03 ;
   RECT 23.18 159.03 157.32 160.74 ;
   RECT 23.18 160.74 157.32 162.45 ;
   RECT 23.18 162.45 157.32 164.16 ;
   RECT 23.18 164.16 157.32 165.87 ;
   RECT 23.18 165.87 157.32 167.58 ;
   RECT 23.18 167.58 157.32 169.29 ;
   RECT 23.18 169.29 157.32 171.0 ;
   RECT 23.18 171.0 157.32 172.71 ;
   RECT 23.18 172.71 157.32 174.42 ;
   RECT 23.18 174.42 157.32 176.13 ;
   RECT 23.18 176.13 157.32 177.84 ;
   RECT 23.18 177.84 157.32 179.55 ;
   RECT 23.18 179.55 157.32 181.26 ;
   RECT 23.18 181.26 157.32 182.97 ;
   RECT 23.18 182.97 157.32 184.68 ;
   RECT 23.18 184.68 157.32 186.39 ;
   RECT 23.18 186.39 157.32 188.1 ;
   RECT 23.18 188.1 157.32 189.81 ;
   RECT 23.18 189.81 157.32 191.52 ;
   RECT 23.18 191.52 157.32 193.23 ;
   RECT 23.18 193.23 157.32 194.94 ;
   RECT 23.18 194.94 157.32 196.65 ;
   RECT 23.18 196.65 157.32 198.36 ;
   RECT 23.18 198.36 157.32 200.07 ;
   RECT 23.18 200.07 157.32 201.78 ;
   RECT 23.18 201.78 157.32 203.49 ;
   RECT 23.18 203.49 157.32 205.2 ;
   RECT 23.18 205.2 157.32 206.91 ;
   RECT 23.18 206.91 157.32 208.62 ;
   RECT 23.18 208.62 157.32 210.33 ;
   RECT 23.18 210.33 157.32 212.04 ;
   RECT 23.18 212.04 157.32 213.75 ;
   RECT 23.18 213.75 157.32 215.46 ;
   RECT 23.18 215.46 157.32 217.17 ;
   RECT 23.18 217.17 157.32 218.88 ;
   RECT 23.18 218.88 157.32 220.59 ;
   RECT 23.18 220.59 157.32 222.3 ;
   RECT 23.18 222.3 157.32 224.01 ;
   RECT 23.18 224.01 157.32 225.72 ;
   RECT 23.18 225.72 157.32 227.43 ;
   RECT 23.18 227.43 157.32 229.14 ;
   RECT 23.18 229.14 157.32 230.85 ;
   RECT 23.18 230.85 157.32 232.56 ;
   RECT 23.18 232.56 157.32 234.27 ;
   RECT 23.18 234.27 157.32 235.98 ;
   RECT 23.18 235.98 157.32 237.69 ;
   RECT 23.18 237.69 157.32 239.4 ;
   RECT 23.18 239.4 157.32 241.11 ;
   RECT 23.18 241.11 157.32 242.82 ;
   RECT 23.18 242.82 157.32 244.53 ;
   RECT 23.18 244.53 157.32 246.24 ;
   RECT 23.18 246.24 157.32 247.95 ;
   RECT 23.18 247.95 157.32 249.66 ;
   RECT 23.18 249.66 157.32 251.37 ;
   RECT 23.18 251.37 157.32 253.08 ;
   RECT 23.18 253.08 157.32 254.79 ;
   RECT 23.18 254.79 157.32 256.5 ;
   RECT 23.18 256.5 157.32 258.21 ;
   RECT 23.18 258.21 157.32 259.92 ;
   RECT 23.18 259.92 157.32 261.63 ;
   RECT 23.18 261.63 157.32 263.34 ;
   RECT 23.18 263.34 157.32 265.05 ;
   RECT 23.18 265.05 157.32 266.76 ;
   RECT 23.18 266.76 157.32 268.47 ;
   RECT 23.18 268.47 157.32 270.18 ;
   RECT 23.18 270.18 157.32 271.89 ;
   RECT 23.18 271.89 157.32 273.6 ;
   RECT 23.18 273.6 157.32 275.31 ;
   RECT 23.18 275.31 157.32 277.02 ;
   RECT 23.18 277.02 157.32 278.73 ;
   RECT 23.18 278.73 157.32 280.44 ;
   RECT 23.18 280.44 157.32 282.15 ;
   RECT 23.18 282.15 157.32 283.86 ;
   RECT 23.18 283.86 157.32 285.57 ;
   RECT 23.18 285.57 157.32 287.28 ;
   RECT 23.18 287.28 157.32 288.99 ;
   RECT 23.18 288.99 157.32 290.7 ;
   RECT 23.18 290.7 157.32 292.41 ;
   RECT 23.18 292.41 157.32 294.12 ;
   RECT 23.18 294.12 157.32 295.83 ;
   RECT 23.18 295.83 157.32 297.54 ;
   RECT 23.18 297.54 157.32 299.25 ;
   RECT 23.18 299.25 157.32 300.96 ;
   RECT 23.18 300.96 157.32 302.67 ;
   RECT 23.18 302.67 157.32 304.38 ;
   RECT 23.18 304.38 157.32 306.09 ;
   RECT 23.18 306.09 157.32 307.8 ;
   RECT 23.18 307.8 157.32 309.51 ;
   RECT 23.18 309.51 157.32 311.22 ;
   RECT 23.18 311.22 157.32 312.93 ;
   RECT 23.18 312.93 157.32 314.64 ;
   RECT 23.18 314.64 157.32 316.35 ;
   RECT 23.18 316.35 157.32 318.06 ;
   RECT 23.18 318.06 157.32 319.77 ;
   RECT 23.18 319.77 157.32 321.48 ;
   RECT 23.18 321.48 157.32 323.19 ;
   RECT 23.18 323.19 157.32 324.9 ;
   RECT 23.18 324.9 157.32 326.61 ;
   RECT 23.18 326.61 157.32 328.32 ;
   RECT 23.18 328.32 157.32 330.03 ;
   RECT 23.18 330.03 157.32 331.74 ;
   RECT 23.18 331.74 157.32 333.45 ;
   RECT 23.18 333.45 157.32 335.16 ;
   RECT 23.18 335.16 157.32 336.87 ;
   RECT 23.18 336.87 157.32 338.58 ;
   RECT 23.18 338.58 157.32 340.29 ;
   RECT 23.18 340.29 157.32 342.0 ;
   RECT 23.18 342.0 157.32 343.71 ;
   RECT 23.18 343.71 157.32 345.42 ;
   RECT 23.18 345.42 157.32 347.13 ;
   RECT 23.18 347.13 157.32 348.84 ;
   RECT 23.18 348.84 157.32 350.55 ;
   RECT 23.18 350.55 157.32 352.26 ;
   RECT 23.18 352.26 157.32 353.97 ;
   RECT 23.18 353.97 157.32 355.68 ;
   RECT 23.18 355.68 157.32 357.39 ;
   RECT 0.0 357.39 157.32 359.1 ;
   RECT 0.0 359.1 157.32 360.81 ;
   RECT 0.0 360.81 157.32 362.52 ;
   RECT 0.0 362.52 157.32 364.23 ;
   RECT 0.0 364.23 157.32 365.94 ;
   RECT 0.0 365.94 157.32 367.65 ;
   RECT 0.0 367.65 157.32 369.36 ;
   RECT 0.0 369.36 157.32 371.07 ;
   RECT 0.0 371.07 157.32 372.78 ;
   RECT 0.0 372.78 157.32 374.49 ;
   RECT 0.0 374.49 157.32 376.2 ;
   RECT 0.0 376.2 157.32 377.91 ;
   RECT 0.0 377.91 157.32 379.62 ;
   RECT 0.0 379.62 157.32 381.33 ;
   RECT 0.0 381.33 157.32 383.04 ;
   RECT 0.0 383.04 157.32 384.75 ;
   RECT 0.0 384.75 157.32 386.46 ;
   RECT 23.18 386.46 157.32 388.17 ;
   RECT 23.18 388.17 157.32 389.88 ;
   RECT 23.18 389.88 157.32 391.59 ;
   RECT 23.18 391.59 157.32 393.3 ;
   RECT 23.18 393.3 157.32 395.01 ;
   RECT 23.18 395.01 157.32 396.72 ;
   RECT 23.18 396.72 157.32 398.43 ;
   RECT 23.18 398.43 157.32 400.14 ;
   RECT 23.18 400.14 157.32 401.85 ;
   RECT 23.18 401.85 157.32 403.56 ;
   RECT 23.18 403.56 157.32 405.27 ;
   RECT 23.18 405.27 157.32 406.98 ;
   RECT 23.18 406.98 157.32 408.69 ;
   RECT 23.18 408.69 157.32 410.4 ;
   RECT 23.18 410.4 157.32 412.11 ;
   RECT 23.18 412.11 157.32 413.82 ;
   RECT 23.18 413.82 157.32 415.53 ;
   RECT 23.18 415.53 157.32 417.24 ;
   RECT 23.18 417.24 157.32 418.95 ;
   RECT 23.18 418.95 157.32 420.66 ;
   RECT 23.18 420.66 157.32 422.37 ;
   RECT 23.18 422.37 157.32 424.08 ;
   RECT 23.18 424.08 157.32 425.79 ;
   RECT 23.18 425.79 157.32 427.5 ;
   RECT 23.18 427.5 157.32 429.21 ;
   RECT 23.18 429.21 157.32 430.92 ;
   RECT 23.18 430.92 157.32 432.63 ;
   RECT 23.18 432.63 157.32 434.34 ;
   RECT 23.18 434.34 157.32 436.05 ;
   RECT 23.18 436.05 157.32 437.76 ;
   RECT 23.18 437.76 157.32 439.47 ;
   RECT 23.18 439.47 157.32 441.18 ;
   RECT 23.18 441.18 157.32 442.89 ;
   RECT 23.18 442.89 157.32 444.6 ;
   RECT 23.18 444.6 157.32 446.31 ;
   RECT 23.18 446.31 157.32 448.02 ;
   RECT 23.18 448.02 157.32 449.73 ;
   RECT 23.18 449.73 157.32 451.44 ;
   RECT 23.18 451.44 157.32 453.15 ;
   RECT 23.18 453.15 157.32 454.86 ;
   RECT 23.18 454.86 157.32 456.57 ;
   RECT 23.18 456.57 157.32 458.28 ;
   RECT 23.18 458.28 157.32 459.99 ;
   RECT 23.18 459.99 157.32 461.7 ;
   RECT 23.18 461.7 157.32 463.41 ;
   RECT 23.18 463.41 157.32 465.12 ;
   RECT 23.18 465.12 157.32 466.83 ;
   RECT 23.18 466.83 157.32 468.54 ;
   RECT 23.18 468.54 157.32 470.25 ;
   RECT 23.18 470.25 157.32 471.96 ;
   RECT 23.18 471.96 157.32 473.67 ;
   RECT 23.18 473.67 157.32 475.38 ;
   RECT 23.18 475.38 157.32 477.09 ;
   RECT 23.18 477.09 157.32 478.8 ;
   RECT 23.18 478.8 157.32 480.51 ;
   RECT 23.18 480.51 157.32 482.22 ;
   RECT 23.18 482.22 157.32 483.93 ;
   RECT 23.18 483.93 157.32 485.64 ;
   RECT 23.18 485.64 157.32 487.35 ;
   RECT 23.18 487.35 157.32 489.06 ;
   RECT 23.18 489.06 157.32 490.77 ;
   RECT 23.18 490.77 157.32 492.48 ;
   RECT 23.18 492.48 157.32 494.19 ;
   RECT 23.18 494.19 157.32 495.9 ;
   RECT 23.18 495.9 157.32 497.61 ;
   RECT 23.18 497.61 157.32 499.32 ;
   RECT 23.18 499.32 157.32 501.03 ;
   RECT 23.18 501.03 157.32 502.74 ;
   RECT 23.18 502.74 157.32 504.45 ;
   RECT 23.18 504.45 157.32 506.16 ;
   RECT 23.18 506.16 157.32 507.87 ;
   RECT 23.18 507.87 157.32 509.58 ;
   RECT 23.18 509.58 157.32 511.29 ;
   RECT 23.18 511.29 157.32 513.0 ;
   RECT 23.18 513.0 157.32 514.71 ;
   RECT 23.18 514.71 157.32 516.42 ;
   RECT 23.18 516.42 157.32 518.13 ;
   RECT 23.18 518.13 157.32 519.84 ;
   RECT 23.18 519.84 157.32 521.55 ;
   RECT 23.18 521.55 157.32 523.26 ;
   RECT 23.18 523.26 157.32 524.97 ;
   RECT 23.18 524.97 157.32 526.68 ;
   RECT 23.18 526.68 157.32 528.39 ;
   RECT 23.18 528.39 157.32 530.1 ;
   RECT 23.18 530.1 157.32 531.81 ;
   RECT 23.18 531.81 157.32 533.52 ;
   RECT 23.18 533.52 157.32 535.23 ;
   RECT 23.18 535.23 157.32 536.94 ;
   RECT 23.18 536.94 157.32 538.65 ;
   RECT 23.18 538.65 157.32 540.36 ;
   RECT 23.18 540.36 157.32 542.07 ;
   RECT 23.18 542.07 157.32 543.78 ;
   RECT 23.18 543.78 157.32 545.49 ;
   RECT 23.18 545.49 157.32 547.2 ;
   RECT 23.18 547.2 157.32 548.91 ;
   RECT 23.18 548.91 157.32 550.62 ;
   RECT 23.18 550.62 157.32 552.33 ;
   RECT 23.18 552.33 157.32 554.04 ;
   RECT 23.18 554.04 157.32 555.75 ;
   RECT 23.18 555.75 157.32 557.46 ;
   RECT 23.18 557.46 157.32 559.17 ;
   RECT 23.18 559.17 157.32 560.88 ;
   RECT 23.18 560.88 157.32 562.59 ;
   RECT 23.18 562.59 157.32 564.3 ;
   RECT 23.18 564.3 157.32 566.01 ;
   RECT 23.18 566.01 157.32 567.72 ;
   RECT 23.18 567.72 157.32 569.43 ;
   RECT 23.18 569.43 157.32 571.14 ;
   RECT 23.18 571.14 157.32 572.85 ;
   RECT 23.18 572.85 157.32 574.56 ;
   RECT 23.18 574.56 157.32 576.27 ;
   RECT 23.18 576.27 157.32 577.98 ;
   RECT 23.18 577.98 157.32 579.69 ;
   RECT 23.18 579.69 157.32 581.4 ;
   RECT 23.18 581.4 157.32 583.11 ;
   RECT 23.18 583.11 157.32 584.82 ;
   RECT 23.18 584.82 157.32 586.53 ;
   RECT 23.18 586.53 157.32 588.24 ;
   RECT 23.18 588.24 157.32 589.95 ;
   RECT 23.18 589.95 157.32 591.66 ;
   RECT 23.18 591.66 157.32 593.37 ;
   RECT 23.18 593.37 157.32 595.08 ;
   RECT 23.18 595.08 157.32 596.79 ;
   RECT 23.18 596.79 157.32 598.5 ;
   RECT 23.18 598.5 157.32 600.21 ;
   RECT 23.18 600.21 157.32 601.92 ;
   RECT 23.18 601.92 157.32 603.63 ;
   RECT 23.18 603.63 157.32 605.34 ;
   RECT 23.18 605.34 157.32 607.05 ;
   RECT 23.18 607.05 157.32 608.76 ;
   RECT 23.18 608.76 157.32 610.47 ;
   RECT 23.18 610.47 157.32 612.18 ;
   RECT 23.18 612.18 157.32 613.89 ;
   RECT 23.18 613.89 157.32 615.6 ;
   RECT 23.18 615.6 157.32 617.31 ;
   RECT 23.18 617.31 157.32 619.02 ;
   RECT 23.18 619.02 157.32 620.73 ;
   RECT 23.18 620.73 157.32 622.44 ;
   RECT 23.18 622.44 157.32 624.15 ;
   RECT 23.18 624.15 157.32 625.86 ;
   RECT 23.18 625.86 157.32 627.57 ;
   RECT 23.18 627.57 157.32 629.28 ;
   RECT 23.18 629.28 157.32 630.99 ;
   RECT 23.18 630.99 157.32 632.7 ;
   RECT 23.18 632.7 157.32 634.41 ;
   RECT 23.18 634.41 157.32 636.12 ;
   RECT 23.18 636.12 157.32 637.83 ;
   RECT 23.18 637.83 157.32 639.54 ;
   RECT 23.18 639.54 157.32 641.25 ;
   RECT 23.18 641.25 157.32 642.96 ;
   RECT 23.18 642.96 157.32 644.67 ;
   RECT 23.18 644.67 157.32 646.38 ;
   RECT 23.18 646.38 157.32 648.09 ;
   RECT 23.18 648.09 157.32 649.8 ;
   RECT 23.18 649.8 157.32 651.51 ;
   RECT 23.18 651.51 157.32 653.22 ;
   RECT 23.18 653.22 157.32 654.93 ;
   RECT 23.18 654.93 157.32 656.64 ;
   RECT 23.18 656.64 157.32 658.35 ;
   RECT 23.18 658.35 157.32 660.06 ;
   RECT 23.18 660.06 157.32 661.77 ;
   RECT 23.18 661.77 157.32 663.48 ;
   RECT 23.18 663.48 157.32 665.19 ;
   RECT 23.18 665.19 157.32 666.9 ;
   RECT 23.18 666.9 157.32 668.61 ;
   RECT 23.18 668.61 157.32 670.32 ;
   RECT 23.18 670.32 157.32 672.03 ;
   RECT 23.18 672.03 157.32 673.74 ;
   RECT 23.18 673.74 157.32 675.45 ;
   RECT 23.18 675.45 157.32 677.16 ;
   RECT 23.18 677.16 157.32 678.87 ;
   RECT 23.18 678.87 157.32 680.58 ;
   RECT 23.18 680.58 157.32 682.29 ;
   RECT 23.18 682.29 157.32 684.0 ;
   RECT 23.18 684.0 157.32 685.71 ;
   RECT 23.18 685.71 157.32 687.42 ;
   RECT 23.18 687.42 157.32 689.13 ;
   RECT 23.18 689.13 157.32 690.84 ;
   RECT 23.18 690.84 157.32 692.55 ;
   RECT 23.18 692.55 157.32 694.26 ;
   RECT 23.18 694.26 157.32 695.97 ;
   RECT 23.18 695.97 157.32 697.68 ;
   RECT 23.18 697.68 157.32 699.39 ;
   RECT 23.18 699.39 157.32 701.1 ;
   RECT 23.18 701.1 157.32 702.81 ;
   RECT 23.18 702.81 157.32 704.52 ;
   RECT 23.18 704.52 157.32 706.23 ;
   RECT 23.18 706.23 157.32 707.94 ;
   RECT 23.18 707.94 157.32 709.65 ;
   RECT 23.18 709.65 157.32 711.36 ;
   RECT 23.18 711.36 157.32 713.07 ;
   RECT 23.18 713.07 157.32 714.78 ;
   RECT 23.18 714.78 157.32 716.49 ;
   RECT 23.18 716.49 157.32 718.2 ;
   RECT 23.18 718.2 157.32 719.91 ;
   RECT 23.18 719.91 157.32 721.62 ;
   RECT 23.18 721.62 157.32 723.33 ;
   RECT 23.18 723.33 157.32 725.04 ;
   RECT 23.18 725.04 157.32 726.75 ;
   RECT 23.18 726.75 157.32 728.46 ;
   RECT 23.18 728.46 157.32 730.17 ;
   RECT 23.18 730.17 157.32 731.88 ;
   RECT 23.18 731.88 157.32 733.59 ;
   RECT 23.18 733.59 157.32 735.3 ;
   RECT 23.18 735.3 157.32 737.01 ;
   RECT 23.18 737.01 157.32 738.72 ;
   RECT 23.18 738.72 157.32 740.43 ;
   RECT 23.18 740.43 157.32 742.14 ;
   RECT 23.18 742.14 157.32 743.85 ;
   RECT 23.18 743.85 157.32 745.56 ;
   RECT 23.18 745.56 157.32 747.27 ;
   RECT 23.18 747.27 157.32 748.98 ;
   RECT 23.18 748.98 157.32 750.69 ;
   RECT 23.18 750.69 157.32 752.4 ;
   RECT 23.18 752.4 157.32 754.11 ;
   RECT 23.18 754.11 157.32 755.82 ;
  LAYER via3 ;
   RECT 23.18 0.0 157.32 1.71 ;
   RECT 23.18 1.71 157.32 3.42 ;
   RECT 23.18 3.42 157.32 5.13 ;
   RECT 23.18 5.13 157.32 6.84 ;
   RECT 23.18 6.84 157.32 8.55 ;
   RECT 23.18 8.55 157.32 10.26 ;
   RECT 23.18 10.26 157.32 11.97 ;
   RECT 23.18 11.97 157.32 13.68 ;
   RECT 23.18 13.68 157.32 15.39 ;
   RECT 23.18 15.39 157.32 17.1 ;
   RECT 23.18 17.1 157.32 18.81 ;
   RECT 23.18 18.81 157.32 20.52 ;
   RECT 23.18 20.52 157.32 22.23 ;
   RECT 23.18 22.23 157.32 23.94 ;
   RECT 23.18 23.94 157.32 25.65 ;
   RECT 23.18 25.65 157.32 27.36 ;
   RECT 23.18 27.36 157.32 29.07 ;
   RECT 23.18 29.07 157.32 30.78 ;
   RECT 23.18 30.78 157.32 32.49 ;
   RECT 23.18 32.49 157.32 34.2 ;
   RECT 23.18 34.2 157.32 35.91 ;
   RECT 23.18 35.91 157.32 37.62 ;
   RECT 23.18 37.62 157.32 39.33 ;
   RECT 23.18 39.33 157.32 41.04 ;
   RECT 23.18 41.04 157.32 42.75 ;
   RECT 23.18 42.75 157.32 44.46 ;
   RECT 23.18 44.46 157.32 46.17 ;
   RECT 23.18 46.17 157.32 47.88 ;
   RECT 23.18 47.88 157.32 49.59 ;
   RECT 23.18 49.59 157.32 51.3 ;
   RECT 23.18 51.3 157.32 53.01 ;
   RECT 23.18 53.01 157.32 54.72 ;
   RECT 23.18 54.72 157.32 56.43 ;
   RECT 23.18 56.43 157.32 58.14 ;
   RECT 23.18 58.14 157.32 59.85 ;
   RECT 23.18 59.85 157.32 61.56 ;
   RECT 23.18 61.56 157.32 63.27 ;
   RECT 23.18 63.27 157.32 64.98 ;
   RECT 23.18 64.98 157.32 66.69 ;
   RECT 23.18 66.69 157.32 68.4 ;
   RECT 23.18 68.4 157.32 70.11 ;
   RECT 23.18 70.11 157.32 71.82 ;
   RECT 23.18 71.82 157.32 73.53 ;
   RECT 23.18 73.53 157.32 75.24 ;
   RECT 23.18 75.24 157.32 76.95 ;
   RECT 23.18 76.95 157.32 78.66 ;
   RECT 23.18 78.66 157.32 80.37 ;
   RECT 23.18 80.37 157.32 82.08 ;
   RECT 23.18 82.08 157.32 83.79 ;
   RECT 23.18 83.79 157.32 85.5 ;
   RECT 23.18 85.5 157.32 87.21 ;
   RECT 23.18 87.21 157.32 88.92 ;
   RECT 23.18 88.92 157.32 90.63 ;
   RECT 23.18 90.63 157.32 92.34 ;
   RECT 23.18 92.34 157.32 94.05 ;
   RECT 23.18 94.05 157.32 95.76 ;
   RECT 23.18 95.76 157.32 97.47 ;
   RECT 23.18 97.47 157.32 99.18 ;
   RECT 23.18 99.18 157.32 100.89 ;
   RECT 23.18 100.89 157.32 102.6 ;
   RECT 23.18 102.6 157.32 104.31 ;
   RECT 23.18 104.31 157.32 106.02 ;
   RECT 23.18 106.02 157.32 107.73 ;
   RECT 23.18 107.73 157.32 109.44 ;
   RECT 23.18 109.44 157.32 111.15 ;
   RECT 23.18 111.15 157.32 112.86 ;
   RECT 23.18 112.86 157.32 114.57 ;
   RECT 23.18 114.57 157.32 116.28 ;
   RECT 23.18 116.28 157.32 117.99 ;
   RECT 23.18 117.99 157.32 119.7 ;
   RECT 23.18 119.7 157.32 121.41 ;
   RECT 23.18 121.41 157.32 123.12 ;
   RECT 23.18 123.12 157.32 124.83 ;
   RECT 23.18 124.83 157.32 126.54 ;
   RECT 23.18 126.54 157.32 128.25 ;
   RECT 23.18 128.25 157.32 129.96 ;
   RECT 23.18 129.96 157.32 131.67 ;
   RECT 23.18 131.67 157.32 133.38 ;
   RECT 23.18 133.38 157.32 135.09 ;
   RECT 23.18 135.09 157.32 136.8 ;
   RECT 23.18 136.8 157.32 138.51 ;
   RECT 23.18 138.51 157.32 140.22 ;
   RECT 23.18 140.22 157.32 141.93 ;
   RECT 23.18 141.93 157.32 143.64 ;
   RECT 23.18 143.64 157.32 145.35 ;
   RECT 23.18 145.35 157.32 147.06 ;
   RECT 23.18 147.06 157.32 148.77 ;
   RECT 23.18 148.77 157.32 150.48 ;
   RECT 23.18 150.48 157.32 152.19 ;
   RECT 23.18 152.19 157.32 153.9 ;
   RECT 23.18 153.9 157.32 155.61 ;
   RECT 23.18 155.61 157.32 157.32 ;
   RECT 23.18 157.32 157.32 159.03 ;
   RECT 23.18 159.03 157.32 160.74 ;
   RECT 23.18 160.74 157.32 162.45 ;
   RECT 23.18 162.45 157.32 164.16 ;
   RECT 23.18 164.16 157.32 165.87 ;
   RECT 23.18 165.87 157.32 167.58 ;
   RECT 23.18 167.58 157.32 169.29 ;
   RECT 23.18 169.29 157.32 171.0 ;
   RECT 23.18 171.0 157.32 172.71 ;
   RECT 23.18 172.71 157.32 174.42 ;
   RECT 23.18 174.42 157.32 176.13 ;
   RECT 23.18 176.13 157.32 177.84 ;
   RECT 23.18 177.84 157.32 179.55 ;
   RECT 23.18 179.55 157.32 181.26 ;
   RECT 23.18 181.26 157.32 182.97 ;
   RECT 23.18 182.97 157.32 184.68 ;
   RECT 23.18 184.68 157.32 186.39 ;
   RECT 23.18 186.39 157.32 188.1 ;
   RECT 23.18 188.1 157.32 189.81 ;
   RECT 23.18 189.81 157.32 191.52 ;
   RECT 23.18 191.52 157.32 193.23 ;
   RECT 23.18 193.23 157.32 194.94 ;
   RECT 23.18 194.94 157.32 196.65 ;
   RECT 23.18 196.65 157.32 198.36 ;
   RECT 23.18 198.36 157.32 200.07 ;
   RECT 23.18 200.07 157.32 201.78 ;
   RECT 23.18 201.78 157.32 203.49 ;
   RECT 23.18 203.49 157.32 205.2 ;
   RECT 23.18 205.2 157.32 206.91 ;
   RECT 23.18 206.91 157.32 208.62 ;
   RECT 23.18 208.62 157.32 210.33 ;
   RECT 23.18 210.33 157.32 212.04 ;
   RECT 23.18 212.04 157.32 213.75 ;
   RECT 23.18 213.75 157.32 215.46 ;
   RECT 23.18 215.46 157.32 217.17 ;
   RECT 23.18 217.17 157.32 218.88 ;
   RECT 23.18 218.88 157.32 220.59 ;
   RECT 23.18 220.59 157.32 222.3 ;
   RECT 23.18 222.3 157.32 224.01 ;
   RECT 23.18 224.01 157.32 225.72 ;
   RECT 23.18 225.72 157.32 227.43 ;
   RECT 23.18 227.43 157.32 229.14 ;
   RECT 23.18 229.14 157.32 230.85 ;
   RECT 23.18 230.85 157.32 232.56 ;
   RECT 23.18 232.56 157.32 234.27 ;
   RECT 23.18 234.27 157.32 235.98 ;
   RECT 23.18 235.98 157.32 237.69 ;
   RECT 23.18 237.69 157.32 239.4 ;
   RECT 23.18 239.4 157.32 241.11 ;
   RECT 23.18 241.11 157.32 242.82 ;
   RECT 23.18 242.82 157.32 244.53 ;
   RECT 23.18 244.53 157.32 246.24 ;
   RECT 23.18 246.24 157.32 247.95 ;
   RECT 23.18 247.95 157.32 249.66 ;
   RECT 23.18 249.66 157.32 251.37 ;
   RECT 23.18 251.37 157.32 253.08 ;
   RECT 23.18 253.08 157.32 254.79 ;
   RECT 23.18 254.79 157.32 256.5 ;
   RECT 23.18 256.5 157.32 258.21 ;
   RECT 23.18 258.21 157.32 259.92 ;
   RECT 23.18 259.92 157.32 261.63 ;
   RECT 23.18 261.63 157.32 263.34 ;
   RECT 23.18 263.34 157.32 265.05 ;
   RECT 23.18 265.05 157.32 266.76 ;
   RECT 23.18 266.76 157.32 268.47 ;
   RECT 23.18 268.47 157.32 270.18 ;
   RECT 23.18 270.18 157.32 271.89 ;
   RECT 23.18 271.89 157.32 273.6 ;
   RECT 23.18 273.6 157.32 275.31 ;
   RECT 23.18 275.31 157.32 277.02 ;
   RECT 23.18 277.02 157.32 278.73 ;
   RECT 23.18 278.73 157.32 280.44 ;
   RECT 23.18 280.44 157.32 282.15 ;
   RECT 23.18 282.15 157.32 283.86 ;
   RECT 23.18 283.86 157.32 285.57 ;
   RECT 23.18 285.57 157.32 287.28 ;
   RECT 23.18 287.28 157.32 288.99 ;
   RECT 23.18 288.99 157.32 290.7 ;
   RECT 23.18 290.7 157.32 292.41 ;
   RECT 23.18 292.41 157.32 294.12 ;
   RECT 23.18 294.12 157.32 295.83 ;
   RECT 23.18 295.83 157.32 297.54 ;
   RECT 23.18 297.54 157.32 299.25 ;
   RECT 23.18 299.25 157.32 300.96 ;
   RECT 23.18 300.96 157.32 302.67 ;
   RECT 23.18 302.67 157.32 304.38 ;
   RECT 23.18 304.38 157.32 306.09 ;
   RECT 23.18 306.09 157.32 307.8 ;
   RECT 23.18 307.8 157.32 309.51 ;
   RECT 23.18 309.51 157.32 311.22 ;
   RECT 23.18 311.22 157.32 312.93 ;
   RECT 23.18 312.93 157.32 314.64 ;
   RECT 23.18 314.64 157.32 316.35 ;
   RECT 23.18 316.35 157.32 318.06 ;
   RECT 23.18 318.06 157.32 319.77 ;
   RECT 23.18 319.77 157.32 321.48 ;
   RECT 23.18 321.48 157.32 323.19 ;
   RECT 23.18 323.19 157.32 324.9 ;
   RECT 23.18 324.9 157.32 326.61 ;
   RECT 23.18 326.61 157.32 328.32 ;
   RECT 23.18 328.32 157.32 330.03 ;
   RECT 23.18 330.03 157.32 331.74 ;
   RECT 23.18 331.74 157.32 333.45 ;
   RECT 23.18 333.45 157.32 335.16 ;
   RECT 23.18 335.16 157.32 336.87 ;
   RECT 23.18 336.87 157.32 338.58 ;
   RECT 23.18 338.58 157.32 340.29 ;
   RECT 23.18 340.29 157.32 342.0 ;
   RECT 23.18 342.0 157.32 343.71 ;
   RECT 23.18 343.71 157.32 345.42 ;
   RECT 23.18 345.42 157.32 347.13 ;
   RECT 23.18 347.13 157.32 348.84 ;
   RECT 23.18 348.84 157.32 350.55 ;
   RECT 23.18 350.55 157.32 352.26 ;
   RECT 23.18 352.26 157.32 353.97 ;
   RECT 23.18 353.97 157.32 355.68 ;
   RECT 23.18 355.68 157.32 357.39 ;
   RECT 0.0 357.39 157.32 359.1 ;
   RECT 0.0 359.1 157.32 360.81 ;
   RECT 0.0 360.81 157.32 362.52 ;
   RECT 0.0 362.52 157.32 364.23 ;
   RECT 0.0 364.23 157.32 365.94 ;
   RECT 0.0 365.94 157.32 367.65 ;
   RECT 0.0 367.65 157.32 369.36 ;
   RECT 0.0 369.36 157.32 371.07 ;
   RECT 0.0 371.07 157.32 372.78 ;
   RECT 0.0 372.78 157.32 374.49 ;
   RECT 0.0 374.49 157.32 376.2 ;
   RECT 0.0 376.2 157.32 377.91 ;
   RECT 0.0 377.91 157.32 379.62 ;
   RECT 0.0 379.62 157.32 381.33 ;
   RECT 0.0 381.33 157.32 383.04 ;
   RECT 0.0 383.04 157.32 384.75 ;
   RECT 0.0 384.75 157.32 386.46 ;
   RECT 23.18 386.46 157.32 388.17 ;
   RECT 23.18 388.17 157.32 389.88 ;
   RECT 23.18 389.88 157.32 391.59 ;
   RECT 23.18 391.59 157.32 393.3 ;
   RECT 23.18 393.3 157.32 395.01 ;
   RECT 23.18 395.01 157.32 396.72 ;
   RECT 23.18 396.72 157.32 398.43 ;
   RECT 23.18 398.43 157.32 400.14 ;
   RECT 23.18 400.14 157.32 401.85 ;
   RECT 23.18 401.85 157.32 403.56 ;
   RECT 23.18 403.56 157.32 405.27 ;
   RECT 23.18 405.27 157.32 406.98 ;
   RECT 23.18 406.98 157.32 408.69 ;
   RECT 23.18 408.69 157.32 410.4 ;
   RECT 23.18 410.4 157.32 412.11 ;
   RECT 23.18 412.11 157.32 413.82 ;
   RECT 23.18 413.82 157.32 415.53 ;
   RECT 23.18 415.53 157.32 417.24 ;
   RECT 23.18 417.24 157.32 418.95 ;
   RECT 23.18 418.95 157.32 420.66 ;
   RECT 23.18 420.66 157.32 422.37 ;
   RECT 23.18 422.37 157.32 424.08 ;
   RECT 23.18 424.08 157.32 425.79 ;
   RECT 23.18 425.79 157.32 427.5 ;
   RECT 23.18 427.5 157.32 429.21 ;
   RECT 23.18 429.21 157.32 430.92 ;
   RECT 23.18 430.92 157.32 432.63 ;
   RECT 23.18 432.63 157.32 434.34 ;
   RECT 23.18 434.34 157.32 436.05 ;
   RECT 23.18 436.05 157.32 437.76 ;
   RECT 23.18 437.76 157.32 439.47 ;
   RECT 23.18 439.47 157.32 441.18 ;
   RECT 23.18 441.18 157.32 442.89 ;
   RECT 23.18 442.89 157.32 444.6 ;
   RECT 23.18 444.6 157.32 446.31 ;
   RECT 23.18 446.31 157.32 448.02 ;
   RECT 23.18 448.02 157.32 449.73 ;
   RECT 23.18 449.73 157.32 451.44 ;
   RECT 23.18 451.44 157.32 453.15 ;
   RECT 23.18 453.15 157.32 454.86 ;
   RECT 23.18 454.86 157.32 456.57 ;
   RECT 23.18 456.57 157.32 458.28 ;
   RECT 23.18 458.28 157.32 459.99 ;
   RECT 23.18 459.99 157.32 461.7 ;
   RECT 23.18 461.7 157.32 463.41 ;
   RECT 23.18 463.41 157.32 465.12 ;
   RECT 23.18 465.12 157.32 466.83 ;
   RECT 23.18 466.83 157.32 468.54 ;
   RECT 23.18 468.54 157.32 470.25 ;
   RECT 23.18 470.25 157.32 471.96 ;
   RECT 23.18 471.96 157.32 473.67 ;
   RECT 23.18 473.67 157.32 475.38 ;
   RECT 23.18 475.38 157.32 477.09 ;
   RECT 23.18 477.09 157.32 478.8 ;
   RECT 23.18 478.8 157.32 480.51 ;
   RECT 23.18 480.51 157.32 482.22 ;
   RECT 23.18 482.22 157.32 483.93 ;
   RECT 23.18 483.93 157.32 485.64 ;
   RECT 23.18 485.64 157.32 487.35 ;
   RECT 23.18 487.35 157.32 489.06 ;
   RECT 23.18 489.06 157.32 490.77 ;
   RECT 23.18 490.77 157.32 492.48 ;
   RECT 23.18 492.48 157.32 494.19 ;
   RECT 23.18 494.19 157.32 495.9 ;
   RECT 23.18 495.9 157.32 497.61 ;
   RECT 23.18 497.61 157.32 499.32 ;
   RECT 23.18 499.32 157.32 501.03 ;
   RECT 23.18 501.03 157.32 502.74 ;
   RECT 23.18 502.74 157.32 504.45 ;
   RECT 23.18 504.45 157.32 506.16 ;
   RECT 23.18 506.16 157.32 507.87 ;
   RECT 23.18 507.87 157.32 509.58 ;
   RECT 23.18 509.58 157.32 511.29 ;
   RECT 23.18 511.29 157.32 513.0 ;
   RECT 23.18 513.0 157.32 514.71 ;
   RECT 23.18 514.71 157.32 516.42 ;
   RECT 23.18 516.42 157.32 518.13 ;
   RECT 23.18 518.13 157.32 519.84 ;
   RECT 23.18 519.84 157.32 521.55 ;
   RECT 23.18 521.55 157.32 523.26 ;
   RECT 23.18 523.26 157.32 524.97 ;
   RECT 23.18 524.97 157.32 526.68 ;
   RECT 23.18 526.68 157.32 528.39 ;
   RECT 23.18 528.39 157.32 530.1 ;
   RECT 23.18 530.1 157.32 531.81 ;
   RECT 23.18 531.81 157.32 533.52 ;
   RECT 23.18 533.52 157.32 535.23 ;
   RECT 23.18 535.23 157.32 536.94 ;
   RECT 23.18 536.94 157.32 538.65 ;
   RECT 23.18 538.65 157.32 540.36 ;
   RECT 23.18 540.36 157.32 542.07 ;
   RECT 23.18 542.07 157.32 543.78 ;
   RECT 23.18 543.78 157.32 545.49 ;
   RECT 23.18 545.49 157.32 547.2 ;
   RECT 23.18 547.2 157.32 548.91 ;
   RECT 23.18 548.91 157.32 550.62 ;
   RECT 23.18 550.62 157.32 552.33 ;
   RECT 23.18 552.33 157.32 554.04 ;
   RECT 23.18 554.04 157.32 555.75 ;
   RECT 23.18 555.75 157.32 557.46 ;
   RECT 23.18 557.46 157.32 559.17 ;
   RECT 23.18 559.17 157.32 560.88 ;
   RECT 23.18 560.88 157.32 562.59 ;
   RECT 23.18 562.59 157.32 564.3 ;
   RECT 23.18 564.3 157.32 566.01 ;
   RECT 23.18 566.01 157.32 567.72 ;
   RECT 23.18 567.72 157.32 569.43 ;
   RECT 23.18 569.43 157.32 571.14 ;
   RECT 23.18 571.14 157.32 572.85 ;
   RECT 23.18 572.85 157.32 574.56 ;
   RECT 23.18 574.56 157.32 576.27 ;
   RECT 23.18 576.27 157.32 577.98 ;
   RECT 23.18 577.98 157.32 579.69 ;
   RECT 23.18 579.69 157.32 581.4 ;
   RECT 23.18 581.4 157.32 583.11 ;
   RECT 23.18 583.11 157.32 584.82 ;
   RECT 23.18 584.82 157.32 586.53 ;
   RECT 23.18 586.53 157.32 588.24 ;
   RECT 23.18 588.24 157.32 589.95 ;
   RECT 23.18 589.95 157.32 591.66 ;
   RECT 23.18 591.66 157.32 593.37 ;
   RECT 23.18 593.37 157.32 595.08 ;
   RECT 23.18 595.08 157.32 596.79 ;
   RECT 23.18 596.79 157.32 598.5 ;
   RECT 23.18 598.5 157.32 600.21 ;
   RECT 23.18 600.21 157.32 601.92 ;
   RECT 23.18 601.92 157.32 603.63 ;
   RECT 23.18 603.63 157.32 605.34 ;
   RECT 23.18 605.34 157.32 607.05 ;
   RECT 23.18 607.05 157.32 608.76 ;
   RECT 23.18 608.76 157.32 610.47 ;
   RECT 23.18 610.47 157.32 612.18 ;
   RECT 23.18 612.18 157.32 613.89 ;
   RECT 23.18 613.89 157.32 615.6 ;
   RECT 23.18 615.6 157.32 617.31 ;
   RECT 23.18 617.31 157.32 619.02 ;
   RECT 23.18 619.02 157.32 620.73 ;
   RECT 23.18 620.73 157.32 622.44 ;
   RECT 23.18 622.44 157.32 624.15 ;
   RECT 23.18 624.15 157.32 625.86 ;
   RECT 23.18 625.86 157.32 627.57 ;
   RECT 23.18 627.57 157.32 629.28 ;
   RECT 23.18 629.28 157.32 630.99 ;
   RECT 23.18 630.99 157.32 632.7 ;
   RECT 23.18 632.7 157.32 634.41 ;
   RECT 23.18 634.41 157.32 636.12 ;
   RECT 23.18 636.12 157.32 637.83 ;
   RECT 23.18 637.83 157.32 639.54 ;
   RECT 23.18 639.54 157.32 641.25 ;
   RECT 23.18 641.25 157.32 642.96 ;
   RECT 23.18 642.96 157.32 644.67 ;
   RECT 23.18 644.67 157.32 646.38 ;
   RECT 23.18 646.38 157.32 648.09 ;
   RECT 23.18 648.09 157.32 649.8 ;
   RECT 23.18 649.8 157.32 651.51 ;
   RECT 23.18 651.51 157.32 653.22 ;
   RECT 23.18 653.22 157.32 654.93 ;
   RECT 23.18 654.93 157.32 656.64 ;
   RECT 23.18 656.64 157.32 658.35 ;
   RECT 23.18 658.35 157.32 660.06 ;
   RECT 23.18 660.06 157.32 661.77 ;
   RECT 23.18 661.77 157.32 663.48 ;
   RECT 23.18 663.48 157.32 665.19 ;
   RECT 23.18 665.19 157.32 666.9 ;
   RECT 23.18 666.9 157.32 668.61 ;
   RECT 23.18 668.61 157.32 670.32 ;
   RECT 23.18 670.32 157.32 672.03 ;
   RECT 23.18 672.03 157.32 673.74 ;
   RECT 23.18 673.74 157.32 675.45 ;
   RECT 23.18 675.45 157.32 677.16 ;
   RECT 23.18 677.16 157.32 678.87 ;
   RECT 23.18 678.87 157.32 680.58 ;
   RECT 23.18 680.58 157.32 682.29 ;
   RECT 23.18 682.29 157.32 684.0 ;
   RECT 23.18 684.0 157.32 685.71 ;
   RECT 23.18 685.71 157.32 687.42 ;
   RECT 23.18 687.42 157.32 689.13 ;
   RECT 23.18 689.13 157.32 690.84 ;
   RECT 23.18 690.84 157.32 692.55 ;
   RECT 23.18 692.55 157.32 694.26 ;
   RECT 23.18 694.26 157.32 695.97 ;
   RECT 23.18 695.97 157.32 697.68 ;
   RECT 23.18 697.68 157.32 699.39 ;
   RECT 23.18 699.39 157.32 701.1 ;
   RECT 23.18 701.1 157.32 702.81 ;
   RECT 23.18 702.81 157.32 704.52 ;
   RECT 23.18 704.52 157.32 706.23 ;
   RECT 23.18 706.23 157.32 707.94 ;
   RECT 23.18 707.94 157.32 709.65 ;
   RECT 23.18 709.65 157.32 711.36 ;
   RECT 23.18 711.36 157.32 713.07 ;
   RECT 23.18 713.07 157.32 714.78 ;
   RECT 23.18 714.78 157.32 716.49 ;
   RECT 23.18 716.49 157.32 718.2 ;
   RECT 23.18 718.2 157.32 719.91 ;
   RECT 23.18 719.91 157.32 721.62 ;
   RECT 23.18 721.62 157.32 723.33 ;
   RECT 23.18 723.33 157.32 725.04 ;
   RECT 23.18 725.04 157.32 726.75 ;
   RECT 23.18 726.75 157.32 728.46 ;
   RECT 23.18 728.46 157.32 730.17 ;
   RECT 23.18 730.17 157.32 731.88 ;
   RECT 23.18 731.88 157.32 733.59 ;
   RECT 23.18 733.59 157.32 735.3 ;
   RECT 23.18 735.3 157.32 737.01 ;
   RECT 23.18 737.01 157.32 738.72 ;
   RECT 23.18 738.72 157.32 740.43 ;
   RECT 23.18 740.43 157.32 742.14 ;
   RECT 23.18 742.14 157.32 743.85 ;
   RECT 23.18 743.85 157.32 745.56 ;
   RECT 23.18 745.56 157.32 747.27 ;
   RECT 23.18 747.27 157.32 748.98 ;
   RECT 23.18 748.98 157.32 750.69 ;
   RECT 23.18 750.69 157.32 752.4 ;
   RECT 23.18 752.4 157.32 754.11 ;
   RECT 23.18 754.11 157.32 755.82 ;
  LAYER metal4 ;
   RECT 23.18 0.0 157.32 1.71 ;
   RECT 23.18 1.71 157.32 3.42 ;
   RECT 23.18 3.42 157.32 5.13 ;
   RECT 23.18 5.13 157.32 6.84 ;
   RECT 23.18 6.84 157.32 8.55 ;
   RECT 23.18 8.55 157.32 10.26 ;
   RECT 23.18 10.26 157.32 11.97 ;
   RECT 23.18 11.97 157.32 13.68 ;
   RECT 23.18 13.68 157.32 15.39 ;
   RECT 23.18 15.39 157.32 17.1 ;
   RECT 23.18 17.1 157.32 18.81 ;
   RECT 23.18 18.81 157.32 20.52 ;
   RECT 23.18 20.52 157.32 22.23 ;
   RECT 23.18 22.23 157.32 23.94 ;
   RECT 23.18 23.94 157.32 25.65 ;
   RECT 23.18 25.65 157.32 27.36 ;
   RECT 23.18 27.36 157.32 29.07 ;
   RECT 23.18 29.07 157.32 30.78 ;
   RECT 23.18 30.78 157.32 32.49 ;
   RECT 23.18 32.49 157.32 34.2 ;
   RECT 23.18 34.2 157.32 35.91 ;
   RECT 23.18 35.91 157.32 37.62 ;
   RECT 23.18 37.62 157.32 39.33 ;
   RECT 23.18 39.33 157.32 41.04 ;
   RECT 23.18 41.04 157.32 42.75 ;
   RECT 23.18 42.75 157.32 44.46 ;
   RECT 23.18 44.46 157.32 46.17 ;
   RECT 23.18 46.17 157.32 47.88 ;
   RECT 23.18 47.88 157.32 49.59 ;
   RECT 23.18 49.59 157.32 51.3 ;
   RECT 23.18 51.3 157.32 53.01 ;
   RECT 23.18 53.01 157.32 54.72 ;
   RECT 23.18 54.72 157.32 56.43 ;
   RECT 23.18 56.43 157.32 58.14 ;
   RECT 23.18 58.14 157.32 59.85 ;
   RECT 23.18 59.85 157.32 61.56 ;
   RECT 23.18 61.56 157.32 63.27 ;
   RECT 23.18 63.27 157.32 64.98 ;
   RECT 23.18 64.98 157.32 66.69 ;
   RECT 23.18 66.69 157.32 68.4 ;
   RECT 23.18 68.4 157.32 70.11 ;
   RECT 23.18 70.11 157.32 71.82 ;
   RECT 23.18 71.82 157.32 73.53 ;
   RECT 23.18 73.53 157.32 75.24 ;
   RECT 23.18 75.24 157.32 76.95 ;
   RECT 23.18 76.95 157.32 78.66 ;
   RECT 23.18 78.66 157.32 80.37 ;
   RECT 23.18 80.37 157.32 82.08 ;
   RECT 23.18 82.08 157.32 83.79 ;
   RECT 23.18 83.79 157.32 85.5 ;
   RECT 23.18 85.5 157.32 87.21 ;
   RECT 23.18 87.21 157.32 88.92 ;
   RECT 23.18 88.92 157.32 90.63 ;
   RECT 23.18 90.63 157.32 92.34 ;
   RECT 23.18 92.34 157.32 94.05 ;
   RECT 23.18 94.05 157.32 95.76 ;
   RECT 23.18 95.76 157.32 97.47 ;
   RECT 23.18 97.47 157.32 99.18 ;
   RECT 23.18 99.18 157.32 100.89 ;
   RECT 23.18 100.89 157.32 102.6 ;
   RECT 23.18 102.6 157.32 104.31 ;
   RECT 23.18 104.31 157.32 106.02 ;
   RECT 23.18 106.02 157.32 107.73 ;
   RECT 23.18 107.73 157.32 109.44 ;
   RECT 23.18 109.44 157.32 111.15 ;
   RECT 23.18 111.15 157.32 112.86 ;
   RECT 23.18 112.86 157.32 114.57 ;
   RECT 23.18 114.57 157.32 116.28 ;
   RECT 23.18 116.28 157.32 117.99 ;
   RECT 23.18 117.99 157.32 119.7 ;
   RECT 23.18 119.7 157.32 121.41 ;
   RECT 23.18 121.41 157.32 123.12 ;
   RECT 23.18 123.12 157.32 124.83 ;
   RECT 23.18 124.83 157.32 126.54 ;
   RECT 23.18 126.54 157.32 128.25 ;
   RECT 23.18 128.25 157.32 129.96 ;
   RECT 23.18 129.96 157.32 131.67 ;
   RECT 23.18 131.67 157.32 133.38 ;
   RECT 23.18 133.38 157.32 135.09 ;
   RECT 23.18 135.09 157.32 136.8 ;
   RECT 23.18 136.8 157.32 138.51 ;
   RECT 23.18 138.51 157.32 140.22 ;
   RECT 23.18 140.22 157.32 141.93 ;
   RECT 23.18 141.93 157.32 143.64 ;
   RECT 23.18 143.64 157.32 145.35 ;
   RECT 23.18 145.35 157.32 147.06 ;
   RECT 23.18 147.06 157.32 148.77 ;
   RECT 23.18 148.77 157.32 150.48 ;
   RECT 23.18 150.48 157.32 152.19 ;
   RECT 23.18 152.19 157.32 153.9 ;
   RECT 23.18 153.9 157.32 155.61 ;
   RECT 23.18 155.61 157.32 157.32 ;
   RECT 23.18 157.32 157.32 159.03 ;
   RECT 23.18 159.03 157.32 160.74 ;
   RECT 23.18 160.74 157.32 162.45 ;
   RECT 23.18 162.45 157.32 164.16 ;
   RECT 23.18 164.16 157.32 165.87 ;
   RECT 23.18 165.87 157.32 167.58 ;
   RECT 23.18 167.58 157.32 169.29 ;
   RECT 23.18 169.29 157.32 171.0 ;
   RECT 23.18 171.0 157.32 172.71 ;
   RECT 23.18 172.71 157.32 174.42 ;
   RECT 23.18 174.42 157.32 176.13 ;
   RECT 23.18 176.13 157.32 177.84 ;
   RECT 23.18 177.84 157.32 179.55 ;
   RECT 23.18 179.55 157.32 181.26 ;
   RECT 23.18 181.26 157.32 182.97 ;
   RECT 23.18 182.97 157.32 184.68 ;
   RECT 23.18 184.68 157.32 186.39 ;
   RECT 23.18 186.39 157.32 188.1 ;
   RECT 23.18 188.1 157.32 189.81 ;
   RECT 23.18 189.81 157.32 191.52 ;
   RECT 23.18 191.52 157.32 193.23 ;
   RECT 23.18 193.23 157.32 194.94 ;
   RECT 23.18 194.94 157.32 196.65 ;
   RECT 23.18 196.65 157.32 198.36 ;
   RECT 23.18 198.36 157.32 200.07 ;
   RECT 23.18 200.07 157.32 201.78 ;
   RECT 23.18 201.78 157.32 203.49 ;
   RECT 23.18 203.49 157.32 205.2 ;
   RECT 23.18 205.2 157.32 206.91 ;
   RECT 23.18 206.91 157.32 208.62 ;
   RECT 23.18 208.62 157.32 210.33 ;
   RECT 23.18 210.33 157.32 212.04 ;
   RECT 23.18 212.04 157.32 213.75 ;
   RECT 23.18 213.75 157.32 215.46 ;
   RECT 23.18 215.46 157.32 217.17 ;
   RECT 23.18 217.17 157.32 218.88 ;
   RECT 23.18 218.88 157.32 220.59 ;
   RECT 23.18 220.59 157.32 222.3 ;
   RECT 23.18 222.3 157.32 224.01 ;
   RECT 23.18 224.01 157.32 225.72 ;
   RECT 23.18 225.72 157.32 227.43 ;
   RECT 23.18 227.43 157.32 229.14 ;
   RECT 23.18 229.14 157.32 230.85 ;
   RECT 23.18 230.85 157.32 232.56 ;
   RECT 23.18 232.56 157.32 234.27 ;
   RECT 23.18 234.27 157.32 235.98 ;
   RECT 23.18 235.98 157.32 237.69 ;
   RECT 23.18 237.69 157.32 239.4 ;
   RECT 23.18 239.4 157.32 241.11 ;
   RECT 23.18 241.11 157.32 242.82 ;
   RECT 23.18 242.82 157.32 244.53 ;
   RECT 23.18 244.53 157.32 246.24 ;
   RECT 23.18 246.24 157.32 247.95 ;
   RECT 23.18 247.95 157.32 249.66 ;
   RECT 23.18 249.66 157.32 251.37 ;
   RECT 23.18 251.37 157.32 253.08 ;
   RECT 23.18 253.08 157.32 254.79 ;
   RECT 23.18 254.79 157.32 256.5 ;
   RECT 23.18 256.5 157.32 258.21 ;
   RECT 23.18 258.21 157.32 259.92 ;
   RECT 23.18 259.92 157.32 261.63 ;
   RECT 23.18 261.63 157.32 263.34 ;
   RECT 23.18 263.34 157.32 265.05 ;
   RECT 23.18 265.05 157.32 266.76 ;
   RECT 23.18 266.76 157.32 268.47 ;
   RECT 23.18 268.47 157.32 270.18 ;
   RECT 23.18 270.18 157.32 271.89 ;
   RECT 23.18 271.89 157.32 273.6 ;
   RECT 23.18 273.6 157.32 275.31 ;
   RECT 23.18 275.31 157.32 277.02 ;
   RECT 23.18 277.02 157.32 278.73 ;
   RECT 23.18 278.73 157.32 280.44 ;
   RECT 23.18 280.44 157.32 282.15 ;
   RECT 23.18 282.15 157.32 283.86 ;
   RECT 23.18 283.86 157.32 285.57 ;
   RECT 23.18 285.57 157.32 287.28 ;
   RECT 23.18 287.28 157.32 288.99 ;
   RECT 23.18 288.99 157.32 290.7 ;
   RECT 23.18 290.7 157.32 292.41 ;
   RECT 23.18 292.41 157.32 294.12 ;
   RECT 23.18 294.12 157.32 295.83 ;
   RECT 23.18 295.83 157.32 297.54 ;
   RECT 23.18 297.54 157.32 299.25 ;
   RECT 23.18 299.25 157.32 300.96 ;
   RECT 23.18 300.96 157.32 302.67 ;
   RECT 23.18 302.67 157.32 304.38 ;
   RECT 23.18 304.38 157.32 306.09 ;
   RECT 23.18 306.09 157.32 307.8 ;
   RECT 23.18 307.8 157.32 309.51 ;
   RECT 23.18 309.51 157.32 311.22 ;
   RECT 23.18 311.22 157.32 312.93 ;
   RECT 23.18 312.93 157.32 314.64 ;
   RECT 23.18 314.64 157.32 316.35 ;
   RECT 23.18 316.35 157.32 318.06 ;
   RECT 23.18 318.06 157.32 319.77 ;
   RECT 23.18 319.77 157.32 321.48 ;
   RECT 23.18 321.48 157.32 323.19 ;
   RECT 23.18 323.19 157.32 324.9 ;
   RECT 23.18 324.9 157.32 326.61 ;
   RECT 23.18 326.61 157.32 328.32 ;
   RECT 23.18 328.32 157.32 330.03 ;
   RECT 23.18 330.03 157.32 331.74 ;
   RECT 23.18 331.74 157.32 333.45 ;
   RECT 23.18 333.45 157.32 335.16 ;
   RECT 23.18 335.16 157.32 336.87 ;
   RECT 23.18 336.87 157.32 338.58 ;
   RECT 23.18 338.58 157.32 340.29 ;
   RECT 23.18 340.29 157.32 342.0 ;
   RECT 23.18 342.0 157.32 343.71 ;
   RECT 23.18 343.71 157.32 345.42 ;
   RECT 23.18 345.42 157.32 347.13 ;
   RECT 23.18 347.13 157.32 348.84 ;
   RECT 23.18 348.84 157.32 350.55 ;
   RECT 23.18 350.55 157.32 352.26 ;
   RECT 23.18 352.26 157.32 353.97 ;
   RECT 23.18 353.97 157.32 355.68 ;
   RECT 23.18 355.68 157.32 357.39 ;
   RECT 0.0 357.39 157.32 359.1 ;
   RECT 0.0 359.1 157.32 360.81 ;
   RECT 0.0 360.81 157.32 362.52 ;
   RECT 0.0 362.52 157.32 364.23 ;
   RECT 0.0 364.23 157.32 365.94 ;
   RECT 0.0 365.94 157.32 367.65 ;
   RECT 0.0 367.65 157.32 369.36 ;
   RECT 0.0 369.36 157.32 371.07 ;
   RECT 0.0 371.07 157.32 372.78 ;
   RECT 0.0 372.78 157.32 374.49 ;
   RECT 0.0 374.49 157.32 376.2 ;
   RECT 0.0 376.2 157.32 377.91 ;
   RECT 0.0 377.91 157.32 379.62 ;
   RECT 0.0 379.62 157.32 381.33 ;
   RECT 0.0 381.33 157.32 383.04 ;
   RECT 0.0 383.04 157.32 384.75 ;
   RECT 0.0 384.75 157.32 386.46 ;
   RECT 23.18 386.46 157.32 388.17 ;
   RECT 23.18 388.17 157.32 389.88 ;
   RECT 23.18 389.88 157.32 391.59 ;
   RECT 23.18 391.59 157.32 393.3 ;
   RECT 23.18 393.3 157.32 395.01 ;
   RECT 23.18 395.01 157.32 396.72 ;
   RECT 23.18 396.72 157.32 398.43 ;
   RECT 23.18 398.43 157.32 400.14 ;
   RECT 23.18 400.14 157.32 401.85 ;
   RECT 23.18 401.85 157.32 403.56 ;
   RECT 23.18 403.56 157.32 405.27 ;
   RECT 23.18 405.27 157.32 406.98 ;
   RECT 23.18 406.98 157.32 408.69 ;
   RECT 23.18 408.69 157.32 410.4 ;
   RECT 23.18 410.4 157.32 412.11 ;
   RECT 23.18 412.11 157.32 413.82 ;
   RECT 23.18 413.82 157.32 415.53 ;
   RECT 23.18 415.53 157.32 417.24 ;
   RECT 23.18 417.24 157.32 418.95 ;
   RECT 23.18 418.95 157.32 420.66 ;
   RECT 23.18 420.66 157.32 422.37 ;
   RECT 23.18 422.37 157.32 424.08 ;
   RECT 23.18 424.08 157.32 425.79 ;
   RECT 23.18 425.79 157.32 427.5 ;
   RECT 23.18 427.5 157.32 429.21 ;
   RECT 23.18 429.21 157.32 430.92 ;
   RECT 23.18 430.92 157.32 432.63 ;
   RECT 23.18 432.63 157.32 434.34 ;
   RECT 23.18 434.34 157.32 436.05 ;
   RECT 23.18 436.05 157.32 437.76 ;
   RECT 23.18 437.76 157.32 439.47 ;
   RECT 23.18 439.47 157.32 441.18 ;
   RECT 23.18 441.18 157.32 442.89 ;
   RECT 23.18 442.89 157.32 444.6 ;
   RECT 23.18 444.6 157.32 446.31 ;
   RECT 23.18 446.31 157.32 448.02 ;
   RECT 23.18 448.02 157.32 449.73 ;
   RECT 23.18 449.73 157.32 451.44 ;
   RECT 23.18 451.44 157.32 453.15 ;
   RECT 23.18 453.15 157.32 454.86 ;
   RECT 23.18 454.86 157.32 456.57 ;
   RECT 23.18 456.57 157.32 458.28 ;
   RECT 23.18 458.28 157.32 459.99 ;
   RECT 23.18 459.99 157.32 461.7 ;
   RECT 23.18 461.7 157.32 463.41 ;
   RECT 23.18 463.41 157.32 465.12 ;
   RECT 23.18 465.12 157.32 466.83 ;
   RECT 23.18 466.83 157.32 468.54 ;
   RECT 23.18 468.54 157.32 470.25 ;
   RECT 23.18 470.25 157.32 471.96 ;
   RECT 23.18 471.96 157.32 473.67 ;
   RECT 23.18 473.67 157.32 475.38 ;
   RECT 23.18 475.38 157.32 477.09 ;
   RECT 23.18 477.09 157.32 478.8 ;
   RECT 23.18 478.8 157.32 480.51 ;
   RECT 23.18 480.51 157.32 482.22 ;
   RECT 23.18 482.22 157.32 483.93 ;
   RECT 23.18 483.93 157.32 485.64 ;
   RECT 23.18 485.64 157.32 487.35 ;
   RECT 23.18 487.35 157.32 489.06 ;
   RECT 23.18 489.06 157.32 490.77 ;
   RECT 23.18 490.77 157.32 492.48 ;
   RECT 23.18 492.48 157.32 494.19 ;
   RECT 23.18 494.19 157.32 495.9 ;
   RECT 23.18 495.9 157.32 497.61 ;
   RECT 23.18 497.61 157.32 499.32 ;
   RECT 23.18 499.32 157.32 501.03 ;
   RECT 23.18 501.03 157.32 502.74 ;
   RECT 23.18 502.74 157.32 504.45 ;
   RECT 23.18 504.45 157.32 506.16 ;
   RECT 23.18 506.16 157.32 507.87 ;
   RECT 23.18 507.87 157.32 509.58 ;
   RECT 23.18 509.58 157.32 511.29 ;
   RECT 23.18 511.29 157.32 513.0 ;
   RECT 23.18 513.0 157.32 514.71 ;
   RECT 23.18 514.71 157.32 516.42 ;
   RECT 23.18 516.42 157.32 518.13 ;
   RECT 23.18 518.13 157.32 519.84 ;
   RECT 23.18 519.84 157.32 521.55 ;
   RECT 23.18 521.55 157.32 523.26 ;
   RECT 23.18 523.26 157.32 524.97 ;
   RECT 23.18 524.97 157.32 526.68 ;
   RECT 23.18 526.68 157.32 528.39 ;
   RECT 23.18 528.39 157.32 530.1 ;
   RECT 23.18 530.1 157.32 531.81 ;
   RECT 23.18 531.81 157.32 533.52 ;
   RECT 23.18 533.52 157.32 535.23 ;
   RECT 23.18 535.23 157.32 536.94 ;
   RECT 23.18 536.94 157.32 538.65 ;
   RECT 23.18 538.65 157.32 540.36 ;
   RECT 23.18 540.36 157.32 542.07 ;
   RECT 23.18 542.07 157.32 543.78 ;
   RECT 23.18 543.78 157.32 545.49 ;
   RECT 23.18 545.49 157.32 547.2 ;
   RECT 23.18 547.2 157.32 548.91 ;
   RECT 23.18 548.91 157.32 550.62 ;
   RECT 23.18 550.62 157.32 552.33 ;
   RECT 23.18 552.33 157.32 554.04 ;
   RECT 23.18 554.04 157.32 555.75 ;
   RECT 23.18 555.75 157.32 557.46 ;
   RECT 23.18 557.46 157.32 559.17 ;
   RECT 23.18 559.17 157.32 560.88 ;
   RECT 23.18 560.88 157.32 562.59 ;
   RECT 23.18 562.59 157.32 564.3 ;
   RECT 23.18 564.3 157.32 566.01 ;
   RECT 23.18 566.01 157.32 567.72 ;
   RECT 23.18 567.72 157.32 569.43 ;
   RECT 23.18 569.43 157.32 571.14 ;
   RECT 23.18 571.14 157.32 572.85 ;
   RECT 23.18 572.85 157.32 574.56 ;
   RECT 23.18 574.56 157.32 576.27 ;
   RECT 23.18 576.27 157.32 577.98 ;
   RECT 23.18 577.98 157.32 579.69 ;
   RECT 23.18 579.69 157.32 581.4 ;
   RECT 23.18 581.4 157.32 583.11 ;
   RECT 23.18 583.11 157.32 584.82 ;
   RECT 23.18 584.82 157.32 586.53 ;
   RECT 23.18 586.53 157.32 588.24 ;
   RECT 23.18 588.24 157.32 589.95 ;
   RECT 23.18 589.95 157.32 591.66 ;
   RECT 23.18 591.66 157.32 593.37 ;
   RECT 23.18 593.37 157.32 595.08 ;
   RECT 23.18 595.08 157.32 596.79 ;
   RECT 23.18 596.79 157.32 598.5 ;
   RECT 23.18 598.5 157.32 600.21 ;
   RECT 23.18 600.21 157.32 601.92 ;
   RECT 23.18 601.92 157.32 603.63 ;
   RECT 23.18 603.63 157.32 605.34 ;
   RECT 23.18 605.34 157.32 607.05 ;
   RECT 23.18 607.05 157.32 608.76 ;
   RECT 23.18 608.76 157.32 610.47 ;
   RECT 23.18 610.47 157.32 612.18 ;
   RECT 23.18 612.18 157.32 613.89 ;
   RECT 23.18 613.89 157.32 615.6 ;
   RECT 23.18 615.6 157.32 617.31 ;
   RECT 23.18 617.31 157.32 619.02 ;
   RECT 23.18 619.02 157.32 620.73 ;
   RECT 23.18 620.73 157.32 622.44 ;
   RECT 23.18 622.44 157.32 624.15 ;
   RECT 23.18 624.15 157.32 625.86 ;
   RECT 23.18 625.86 157.32 627.57 ;
   RECT 23.18 627.57 157.32 629.28 ;
   RECT 23.18 629.28 157.32 630.99 ;
   RECT 23.18 630.99 157.32 632.7 ;
   RECT 23.18 632.7 157.32 634.41 ;
   RECT 23.18 634.41 157.32 636.12 ;
   RECT 23.18 636.12 157.32 637.83 ;
   RECT 23.18 637.83 157.32 639.54 ;
   RECT 23.18 639.54 157.32 641.25 ;
   RECT 23.18 641.25 157.32 642.96 ;
   RECT 23.18 642.96 157.32 644.67 ;
   RECT 23.18 644.67 157.32 646.38 ;
   RECT 23.18 646.38 157.32 648.09 ;
   RECT 23.18 648.09 157.32 649.8 ;
   RECT 23.18 649.8 157.32 651.51 ;
   RECT 23.18 651.51 157.32 653.22 ;
   RECT 23.18 653.22 157.32 654.93 ;
   RECT 23.18 654.93 157.32 656.64 ;
   RECT 23.18 656.64 157.32 658.35 ;
   RECT 23.18 658.35 157.32 660.06 ;
   RECT 23.18 660.06 157.32 661.77 ;
   RECT 23.18 661.77 157.32 663.48 ;
   RECT 23.18 663.48 157.32 665.19 ;
   RECT 23.18 665.19 157.32 666.9 ;
   RECT 23.18 666.9 157.32 668.61 ;
   RECT 23.18 668.61 157.32 670.32 ;
   RECT 23.18 670.32 157.32 672.03 ;
   RECT 23.18 672.03 157.32 673.74 ;
   RECT 23.18 673.74 157.32 675.45 ;
   RECT 23.18 675.45 157.32 677.16 ;
   RECT 23.18 677.16 157.32 678.87 ;
   RECT 23.18 678.87 157.32 680.58 ;
   RECT 23.18 680.58 157.32 682.29 ;
   RECT 23.18 682.29 157.32 684.0 ;
   RECT 23.18 684.0 157.32 685.71 ;
   RECT 23.18 685.71 157.32 687.42 ;
   RECT 23.18 687.42 157.32 689.13 ;
   RECT 23.18 689.13 157.32 690.84 ;
   RECT 23.18 690.84 157.32 692.55 ;
   RECT 23.18 692.55 157.32 694.26 ;
   RECT 23.18 694.26 157.32 695.97 ;
   RECT 23.18 695.97 157.32 697.68 ;
   RECT 23.18 697.68 157.32 699.39 ;
   RECT 23.18 699.39 157.32 701.1 ;
   RECT 23.18 701.1 157.32 702.81 ;
   RECT 23.18 702.81 157.32 704.52 ;
   RECT 23.18 704.52 157.32 706.23 ;
   RECT 23.18 706.23 157.32 707.94 ;
   RECT 23.18 707.94 157.32 709.65 ;
   RECT 23.18 709.65 157.32 711.36 ;
   RECT 23.18 711.36 157.32 713.07 ;
   RECT 23.18 713.07 157.32 714.78 ;
   RECT 23.18 714.78 157.32 716.49 ;
   RECT 23.18 716.49 157.32 718.2 ;
   RECT 23.18 718.2 157.32 719.91 ;
   RECT 23.18 719.91 157.32 721.62 ;
   RECT 23.18 721.62 157.32 723.33 ;
   RECT 23.18 723.33 157.32 725.04 ;
   RECT 23.18 725.04 157.32 726.75 ;
   RECT 23.18 726.75 157.32 728.46 ;
   RECT 23.18 728.46 157.32 730.17 ;
   RECT 23.18 730.17 157.32 731.88 ;
   RECT 23.18 731.88 157.32 733.59 ;
   RECT 23.18 733.59 157.32 735.3 ;
   RECT 23.18 735.3 157.32 737.01 ;
   RECT 23.18 737.01 157.32 738.72 ;
   RECT 23.18 738.72 157.32 740.43 ;
   RECT 23.18 740.43 157.32 742.14 ;
   RECT 23.18 742.14 157.32 743.85 ;
   RECT 23.18 743.85 157.32 745.56 ;
   RECT 23.18 745.56 157.32 747.27 ;
   RECT 23.18 747.27 157.32 748.98 ;
   RECT 23.18 748.98 157.32 750.69 ;
   RECT 23.18 750.69 157.32 752.4 ;
   RECT 23.18 752.4 157.32 754.11 ;
   RECT 23.18 754.11 157.32 755.82 ;
 END
END block_414x3978_702

MACRO block_416x441_104
 CLASS BLOCK ;
 FOREIGN block_416x441_104 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 158.08 BY 83.79 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 64.315 154.945 64.885 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 74.955 3.325 75.525 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 20.615 154.945 21.185 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 4.655 3.325 5.225 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 8.075 3.325 8.645 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 9.215 3.325 9.785 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 12.635 3.325 13.205 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 24.415 3.325 24.985 ;
  END
 END o7
 PIN o8
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 25.555 3.325 26.125 ;
  END
 END o8
 PIN o9
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 26.315 3.325 26.885 ;
  END
 END o9
 PIN o10
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 27.455 3.325 28.025 ;
  END
 END o10
 PIN o11
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 28.975 3.325 29.545 ;
  END
 END o11
 PIN o12
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 22.895 3.325 23.465 ;
  END
 END o12
 PIN o13
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 32.015 3.325 32.585 ;
  END
 END o13
 PIN o14
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 33.535 3.325 34.105 ;
  END
 END o14
 PIN o15
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 34.295 3.325 34.865 ;
  END
 END o15
 PIN o16
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 35.055 3.325 35.625 ;
  END
 END o16
 PIN o17
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 35.815 3.325 36.385 ;
  END
 END o17
 PIN o18
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 30.875 3.325 31.445 ;
  END
 END o18
 PIN o19
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 38.855 3.325 39.425 ;
  END
 END o19
 PIN o20
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 39.615 3.325 40.185 ;
  END
 END o20
 PIN o21
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 40.375 3.325 40.945 ;
  END
 END o21
 PIN o22
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 41.135 3.325 41.705 ;
  END
 END o22
 PIN o23
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 42.655 3.325 43.225 ;
  END
 END o23
 PIN o24
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 38.095 3.325 38.665 ;
  END
 END o24
 PIN o25
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 44.935 3.325 45.505 ;
  END
 END o25
 PIN o26
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 45.695 3.325 46.265 ;
  END
 END o26
 PIN o27
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 47.215 3.325 47.785 ;
  END
 END o27
 PIN o28
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 47.975 3.325 48.545 ;
  END
 END o28
 PIN o29
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 48.735 3.325 49.305 ;
  END
 END o29
 PIN o30
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 44.175 3.325 44.745 ;
  END
 END o30
 PIN o31
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 51.775 3.325 52.345 ;
  END
 END o31
 PIN o32
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 52.535 3.325 53.105 ;
  END
 END o32
 PIN o33
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 53.295 3.325 53.865 ;
  END
 END o33
 PIN o34
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 54.055 3.325 54.625 ;
  END
 END o34
 PIN o35
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 54.815 3.325 55.385 ;
  END
 END o35
 PIN o36
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 50.255 3.325 50.825 ;
  END
 END o36
 PIN o37
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 57.855 3.325 58.425 ;
  END
 END o37
 PIN o38
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 58.615 3.325 59.185 ;
  END
 END o38
 PIN o39
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 59.375 3.325 59.945 ;
  END
 END o39
 PIN o40
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 60.895 3.325 61.465 ;
  END
 END o40
 PIN o41
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 61.655 3.325 62.225 ;
  END
 END o41
 PIN o42
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 57.095 3.325 57.665 ;
  END
 END o42
 PIN o43
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 63.935 3.325 64.505 ;
  END
 END o43
 PIN o44
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 65.455 3.325 66.025 ;
  END
 END o44
 PIN o45
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 66.215 3.325 66.785 ;
  END
 END o45
 PIN o46
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 66.975 3.325 67.545 ;
  END
 END o46
 PIN o47
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 67.735 3.325 68.305 ;
  END
 END o47
 PIN o48
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 63.175 3.325 63.745 ;
  END
 END o48
 PIN o49
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 70.775 3.325 71.345 ;
  END
 END o49
 PIN o50
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 71.535 3.325 72.105 ;
  END
 END o50
 PIN o51
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 72.295 3.325 72.865 ;
  END
 END o51
 PIN o52
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 72.675 4.085 73.245 ;
  END
 END o52
 PIN o53
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 73.055 3.325 73.625 ;
  END
 END o53
 PIN o54
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 70.015 3.325 70.585 ;
  END
 END o54
 PIN o55
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 24.415 154.945 24.985 ;
  END
 END o55
 PIN o56
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 25.175 154.945 25.745 ;
  END
 END o56
 PIN o57
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 25.935 154.945 26.505 ;
  END
 END o57
 PIN o58
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 22.895 154.945 23.465 ;
  END
 END o58
 PIN o59
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 29.735 154.945 30.305 ;
  END
 END o59
 PIN o60
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 30.495 154.945 31.065 ;
  END
 END o60
 PIN o61
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 31.255 154.945 31.825 ;
  END
 END o61
 PIN o62
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 28.975 154.945 29.545 ;
  END
 END o62
 PIN o63
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 22.135 154.945 22.705 ;
  END
 END o63
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 51.775 154.945 52.345 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 66.975 154.945 67.545 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 49.495 154.945 50.065 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 50.255 154.945 50.825 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 54.055 154.945 54.625 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 53.295 154.945 53.865 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 47.215 154.945 47.785 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 47.975 154.945 48.545 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 3.515 3.325 4.085 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 19.855 154.945 20.425 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 18.335 154.945 18.905 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 17.575 154.945 18.145 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 48.735 154.945 49.305 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 45.695 154.945 46.265 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 44.935 154.945 45.505 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 74.575 4.085 75.145 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 21.375 154.945 21.945 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 57.095 154.945 57.665 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 57.855 154.945 58.425 ;
  END
 END i18
 PIN i19
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 58.615 154.945 59.185 ;
  END
 END i19
 PIN i20
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 59.375 154.945 59.945 ;
  END
 END i20
 PIN i21
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 60.895 154.945 61.465 ;
  END
 END i21
 PIN i22
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 61.655 154.945 62.225 ;
  END
 END i22
 PIN i23
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 62.415 154.945 62.985 ;
  END
 END i23
 PIN i24
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 63.175 154.945 63.745 ;
  END
 END i24
 PIN i25
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 3.135 154.945 3.705 ;
  END
 END i25
 PIN i26
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 3.895 154.945 4.465 ;
  END
 END i26
 PIN i27
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 4.655 154.945 5.225 ;
  END
 END i27
 PIN i28
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 6.175 154.945 6.745 ;
  END
 END i28
 PIN i29
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 6.935 154.945 7.505 ;
  END
 END i29
 PIN i30
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 7.695 154.945 8.265 ;
  END
 END i30
 PIN i31
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 8.455 154.945 9.025 ;
  END
 END i31
 PIN i32
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 9.215 154.945 9.785 ;
  END
 END i32
 PIN i33
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 10.735 154.945 11.305 ;
  END
 END i33
 PIN i34
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 11.495 154.945 12.065 ;
  END
 END i34
 PIN i35
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 12.255 154.945 12.825 ;
  END
 END i35
 PIN i36
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 13.015 154.945 13.585 ;
  END
 END i36
 PIN i37
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 13.775 154.945 14.345 ;
  END
 END i37
 PIN i38
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 15.295 154.945 15.865 ;
  END
 END i38
 PIN i39
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 16.055 154.945 16.625 ;
  END
 END i39
 OBS
  LAYER metal1 ;
   RECT 0 0 158.08 83.79 ;
  LAYER via1 ;
   RECT 0 0 158.08 83.79 ;
  LAYER metal2 ;
   RECT 0 0 158.08 83.79 ;
  LAYER via2 ;
   RECT 0 0 158.08 83.79 ;
  LAYER metal3 ;
   RECT 0 0 158.08 83.79 ;
  LAYER via3 ;
   RECT 0 0 158.08 83.79 ;
  LAYER metal4 ;
   RECT 0 0 158.08 83.79 ;
 END
END block_416x441_104

MACRO block_414x3969_702
 CLASS BLOCK ;
 FOREIGN block_414x3969_702 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 157.32 BY 754.11 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 749.075 26.885 749.645 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 744.895 26.885 745.465 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 708.225 26.885 708.795 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 256.595 26.885 257.165 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 252.415 26.885 252.985 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 248.425 26.885 248.995 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 244.245 26.885 244.815 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 240.255 26.885 240.825 ;
  END
 END o7
 PIN o8
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 236.075 26.885 236.645 ;
  END
 END o8
 PIN o9
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 232.085 26.885 232.655 ;
  END
 END o9
 PIN o10
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 227.905 26.885 228.475 ;
  END
 END o10
 PIN o11
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 223.915 26.885 224.485 ;
  END
 END o11
 PIN o12
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 219.735 26.885 220.305 ;
  END
 END o12
 PIN o13
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 704.045 26.885 704.615 ;
  END
 END o13
 PIN o14
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 215.745 26.885 216.315 ;
  END
 END o14
 PIN o15
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 211.565 26.885 212.135 ;
  END
 END o15
 PIN o16
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 207.575 26.885 208.145 ;
  END
 END o16
 PIN o17
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 203.395 26.885 203.965 ;
  END
 END o17
 PIN o18
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 199.405 26.885 199.975 ;
  END
 END o18
 PIN o19
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 195.225 26.885 195.795 ;
  END
 END o19
 PIN o20
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 191.235 26.885 191.805 ;
  END
 END o20
 PIN o21
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 187.055 26.885 187.625 ;
  END
 END o21
 PIN o22
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 183.065 26.885 183.635 ;
  END
 END o22
 PIN o23
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 173.755 26.885 174.325 ;
  END
 END o23
 PIN o24
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 700.055 26.885 700.625 ;
  END
 END o24
 PIN o25
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 169.765 26.885 170.335 ;
  END
 END o25
 PIN o26
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 165.585 26.885 166.155 ;
  END
 END o26
 PIN o27
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 161.595 26.885 162.165 ;
  END
 END o27
 PIN o28
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 157.415 26.885 157.985 ;
  END
 END o28
 PIN o29
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 153.425 26.885 153.995 ;
  END
 END o29
 PIN o30
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 149.245 26.885 149.815 ;
  END
 END o30
 PIN o31
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 145.255 26.885 145.825 ;
  END
 END o31
 PIN o32
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 141.075 26.885 141.645 ;
  END
 END o32
 PIN o33
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 137.085 26.885 137.655 ;
  END
 END o33
 PIN o34
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 132.905 26.885 133.475 ;
  END
 END o34
 PIN o35
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 695.875 26.885 696.445 ;
  END
 END o35
 PIN o36
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 128.915 26.885 129.485 ;
  END
 END o36
 PIN o37
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 124.735 26.885 125.305 ;
  END
 END o37
 PIN o38
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 120.745 26.885 121.315 ;
  END
 END o38
 PIN o39
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 116.565 26.885 117.135 ;
  END
 END o39
 PIN o40
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 112.575 26.885 113.145 ;
  END
 END o40
 PIN o41
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 108.395 26.885 108.965 ;
  END
 END o41
 PIN o42
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 104.405 26.885 104.975 ;
  END
 END o42
 PIN o43
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 100.225 26.885 100.795 ;
  END
 END o43
 PIN o44
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 77.995 26.885 78.565 ;
  END
 END o44
 PIN o45
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 73.815 26.885 74.385 ;
  END
 END o45
 PIN o46
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 691.885 26.885 692.455 ;
  END
 END o46
 PIN o47
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 69.825 26.885 70.395 ;
  END
 END o47
 PIN o48
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 65.645 26.885 66.215 ;
  END
 END o48
 PIN o49
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 61.655 26.885 62.225 ;
  END
 END o49
 PIN o50
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 57.475 26.885 58.045 ;
  END
 END o50
 PIN o51
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 53.485 26.885 54.055 ;
  END
 END o51
 PIN o52
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 49.305 26.885 49.875 ;
  END
 END o52
 PIN o53
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 45.315 26.885 45.885 ;
  END
 END o53
 PIN o54
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 41.135 26.885 41.705 ;
  END
 END o54
 PIN o55
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 37.145 26.885 37.715 ;
  END
 END o55
 PIN o56
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 32.965 26.885 33.535 ;
  END
 END o56
 PIN o57
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 687.705 26.885 688.275 ;
  END
 END o57
 PIN o58
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 28.975 26.885 29.545 ;
  END
 END o58
 PIN o59
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 24.795 26.885 25.365 ;
  END
 END o59
 PIN o60
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 20.805 26.885 21.375 ;
  END
 END o60
 PIN o61
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 16.625 26.885 17.195 ;
  END
 END o61
 PIN o62
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 12.635 26.885 13.205 ;
  END
 END o62
 PIN o63
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 8.455 26.885 9.025 ;
  END
 END o63
 PIN o64
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 4.465 26.885 5.035 ;
  END
 END o64
 PIN o65
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 683.715 26.885 684.285 ;
  END
 END o65
 PIN o66
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 679.535 26.885 680.105 ;
  END
 END o66
 PIN o67
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 675.545 26.885 676.115 ;
  END
 END o67
 PIN o68
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 671.365 26.885 671.935 ;
  END
 END o68
 PIN o69
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 740.905 26.885 741.475 ;
  END
 END o69
 PIN o70
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 649.135 26.885 649.705 ;
  END
 END o70
 PIN o71
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 644.955 26.885 645.525 ;
  END
 END o71
 PIN o72
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 640.965 26.885 641.535 ;
  END
 END o72
 PIN o73
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 636.785 26.885 637.355 ;
  END
 END o73
 PIN o74
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 632.795 26.885 633.365 ;
  END
 END o74
 PIN o75
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 628.615 26.885 629.185 ;
  END
 END o75
 PIN o76
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 624.625 26.885 625.195 ;
  END
 END o76
 PIN o77
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 620.445 26.885 621.015 ;
  END
 END o77
 PIN o78
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 616.455 26.885 617.025 ;
  END
 END o78
 PIN o79
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 612.275 26.885 612.845 ;
  END
 END o79
 PIN o80
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 736.725 26.885 737.295 ;
  END
 END o80
 PIN o81
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 608.285 26.885 608.855 ;
  END
 END o81
 PIN o82
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 604.105 26.885 604.675 ;
  END
 END o82
 PIN o83
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 600.115 26.885 600.685 ;
  END
 END o83
 PIN o84
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 595.935 26.885 596.505 ;
  END
 END o84
 PIN o85
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 591.945 26.885 592.515 ;
  END
 END o85
 PIN o86
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 587.765 26.885 588.335 ;
  END
 END o86
 PIN o87
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 583.775 26.885 584.345 ;
  END
 END o87
 PIN o88
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 579.595 26.885 580.165 ;
  END
 END o88
 PIN o89
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 575.605 26.885 576.175 ;
  END
 END o89
 PIN o90
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 571.425 26.885 571.995 ;
  END
 END o90
 PIN o91
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 732.735 26.885 733.305 ;
  END
 END o91
 PIN o92
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 562.305 26.885 562.875 ;
  END
 END o92
 PIN o93
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 558.125 26.885 558.695 ;
  END
 END o93
 PIN o94
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 554.135 26.885 554.705 ;
  END
 END o94
 PIN o95
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 549.955 26.885 550.525 ;
  END
 END o95
 PIN o96
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 545.965 26.885 546.535 ;
  END
 END o96
 PIN o97
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 541.785 26.885 542.355 ;
  END
 END o97
 PIN o98
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 537.795 26.885 538.365 ;
  END
 END o98
 PIN o99
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 533.615 26.885 534.185 ;
  END
 END o99
 PIN o100
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 529.625 26.885 530.195 ;
  END
 END o100
 PIN o101
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 525.445 26.885 526.015 ;
  END
 END o101
 PIN o102
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 728.555 26.885 729.125 ;
  END
 END o102
 PIN o103
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 521.455 26.885 522.025 ;
  END
 END o103
 PIN o104
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 517.275 26.885 517.845 ;
  END
 END o104
 PIN o105
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 513.285 26.885 513.855 ;
  END
 END o105
 PIN o106
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 509.105 26.885 509.675 ;
  END
 END o106
 PIN o107
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 505.115 26.885 505.685 ;
  END
 END o107
 PIN o108
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 500.935 26.885 501.505 ;
  END
 END o108
 PIN o109
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 496.945 26.885 497.515 ;
  END
 END o109
 PIN o110
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 492.765 26.885 493.335 ;
  END
 END o110
 PIN o111
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 488.775 26.885 489.345 ;
  END
 END o111
 PIN o112
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 484.595 26.885 485.165 ;
  END
 END o112
 PIN o113
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 724.565 26.885 725.135 ;
  END
 END o113
 PIN o114
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 462.365 26.885 462.935 ;
  END
 END o114
 PIN o115
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 458.185 26.885 458.755 ;
  END
 END o115
 PIN o116
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 454.195 26.885 454.765 ;
  END
 END o116
 PIN o117
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 450.015 26.885 450.585 ;
  END
 END o117
 PIN o118
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 446.025 26.885 446.595 ;
  END
 END o118
 PIN o119
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 441.845 26.885 442.415 ;
  END
 END o119
 PIN o120
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 437.855 26.885 438.425 ;
  END
 END o120
 PIN o121
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 433.675 26.885 434.245 ;
  END
 END o121
 PIN o122
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 429.685 26.885 430.255 ;
  END
 END o122
 PIN o123
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 425.505 26.885 426.075 ;
  END
 END o123
 PIN o124
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 720.385 26.885 720.955 ;
  END
 END o124
 PIN o125
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 421.515 26.885 422.085 ;
  END
 END o125
 PIN o126
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 417.335 26.885 417.905 ;
  END
 END o126
 PIN o127
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 413.345 26.885 413.915 ;
  END
 END o127
 PIN o128
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 409.165 26.885 409.735 ;
  END
 END o128
 PIN o129
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 405.175 26.885 405.745 ;
  END
 END o129
 PIN o130
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 400.995 26.885 401.565 ;
  END
 END o130
 PIN o131
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 397.005 26.885 397.575 ;
  END
 END o131
 PIN o132
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 392.825 26.885 393.395 ;
  END
 END o132
 PIN o133
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 388.835 26.885 389.405 ;
  END
 END o133
 PIN o134
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 384.655 26.885 385.225 ;
  END
 END o134
 PIN o135
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 716.395 26.885 716.965 ;
  END
 END o135
 PIN o136
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 356.535 26.885 357.105 ;
  END
 END o136
 PIN o137
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 352.355 26.885 352.925 ;
  END
 END o137
 PIN o138
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 348.365 26.885 348.935 ;
  END
 END o138
 PIN o139
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 344.185 26.885 344.755 ;
  END
 END o139
 PIN o140
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 340.195 26.885 340.765 ;
  END
 END o140
 PIN o141
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 336.015 26.885 336.585 ;
  END
 END o141
 PIN o142
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 332.025 26.885 332.595 ;
  END
 END o142
 PIN o143
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 327.845 26.885 328.415 ;
  END
 END o143
 PIN o144
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 323.855 26.885 324.425 ;
  END
 END o144
 PIN o145
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 319.675 26.885 320.245 ;
  END
 END o145
 PIN o146
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 712.215 26.885 712.785 ;
  END
 END o146
 PIN o147
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 315.685 26.885 316.255 ;
  END
 END o147
 PIN o148
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 311.505 26.885 312.075 ;
  END
 END o148
 PIN o149
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 307.515 26.885 308.085 ;
  END
 END o149
 PIN o150
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 303.335 26.885 303.905 ;
  END
 END o150
 PIN o151
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 299.345 26.885 299.915 ;
  END
 END o151
 PIN o152
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 295.165 26.885 295.735 ;
  END
 END o152
 PIN o153
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 291.175 26.885 291.745 ;
  END
 END o153
 PIN o154
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 286.995 26.885 287.565 ;
  END
 END o154
 PIN o155
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 283.005 26.885 283.575 ;
  END
 END o155
 PIN o156
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 278.825 26.885 279.395 ;
  END
 END o156
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 381.805 3.705 382.375 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 364.705 3.705 365.275 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 376.485 3.705 377.055 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 381.425 4.465 381.995 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 382.185 4.465 382.755 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 382.565 3.705 383.135 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 372.875 3.705 373.445 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 359.765 3.705 360.335 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 365.465 3.705 366.035 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 363.375 3.705 363.945 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 360.905 3.705 361.475 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 359.385 4.465 359.955 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 13.015 382.945 13.585 383.515 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 13.015 369.645 13.585 370.215 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 750.785 26.885 751.355 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 746.605 26.885 747.175 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 709.935 26.885 710.505 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 254.885 26.885 255.455 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 250.705 26.885 251.275 ;
  END
 END i18
 PIN i19
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 246.715 26.885 247.285 ;
  END
 END i19
 PIN i20
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 242.535 26.885 243.105 ;
  END
 END i20
 PIN i21
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 238.545 26.885 239.115 ;
  END
 END i21
 PIN i22
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 234.365 26.885 234.935 ;
  END
 END i22
 PIN i23
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 230.375 26.885 230.945 ;
  END
 END i23
 PIN i24
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 226.195 26.885 226.765 ;
  END
 END i24
 PIN i25
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 222.205 26.885 222.775 ;
  END
 END i25
 PIN i26
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 218.025 26.885 218.595 ;
  END
 END i26
 PIN i27
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 705.755 26.885 706.325 ;
  END
 END i27
 PIN i28
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 214.035 26.885 214.605 ;
  END
 END i28
 PIN i29
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 209.855 26.885 210.425 ;
  END
 END i29
 PIN i30
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 205.865 26.885 206.435 ;
  END
 END i30
 PIN i31
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 201.685 26.885 202.255 ;
  END
 END i31
 PIN i32
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 197.695 26.885 198.265 ;
  END
 END i32
 PIN i33
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 193.515 26.885 194.085 ;
  END
 END i33
 PIN i34
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 189.525 26.885 190.095 ;
  END
 END i34
 PIN i35
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 185.345 26.885 185.915 ;
  END
 END i35
 PIN i36
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 181.355 26.885 181.925 ;
  END
 END i36
 PIN i37
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 172.045 26.885 172.615 ;
  END
 END i37
 PIN i38
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 701.765 26.885 702.335 ;
  END
 END i38
 PIN i39
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 168.055 26.885 168.625 ;
  END
 END i39
 PIN i40
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 163.875 26.885 164.445 ;
  END
 END i40
 PIN i41
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 159.885 26.885 160.455 ;
  END
 END i41
 PIN i42
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 155.705 26.885 156.275 ;
  END
 END i42
 PIN i43
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 151.715 26.885 152.285 ;
  END
 END i43
 PIN i44
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 147.535 26.885 148.105 ;
  END
 END i44
 PIN i45
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 143.545 26.885 144.115 ;
  END
 END i45
 PIN i46
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 139.365 26.885 139.935 ;
  END
 END i46
 PIN i47
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 135.375 26.885 135.945 ;
  END
 END i47
 PIN i48
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 131.195 26.885 131.765 ;
  END
 END i48
 PIN i49
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 697.585 26.885 698.155 ;
  END
 END i49
 PIN i50
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 127.205 26.885 127.775 ;
  END
 END i50
 PIN i51
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 123.025 26.885 123.595 ;
  END
 END i51
 PIN i52
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 119.035 26.885 119.605 ;
  END
 END i52
 PIN i53
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 114.855 26.885 115.425 ;
  END
 END i53
 PIN i54
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 110.865 26.885 111.435 ;
  END
 END i54
 PIN i55
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 106.685 26.885 107.255 ;
  END
 END i55
 PIN i56
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 102.695 26.885 103.265 ;
  END
 END i56
 PIN i57
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 98.515 26.885 99.085 ;
  END
 END i57
 PIN i58
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 76.285 26.885 76.855 ;
  END
 END i58
 PIN i59
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 72.105 26.885 72.675 ;
  END
 END i59
 PIN i60
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 693.595 26.885 694.165 ;
  END
 END i60
 PIN i61
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 68.115 26.885 68.685 ;
  END
 END i61
 PIN i62
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 63.935 26.885 64.505 ;
  END
 END i62
 PIN i63
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 59.945 26.885 60.515 ;
  END
 END i63
 PIN i64
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 55.765 26.885 56.335 ;
  END
 END i64
 PIN i65
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 51.775 26.885 52.345 ;
  END
 END i65
 PIN i66
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 47.595 26.885 48.165 ;
  END
 END i66
 PIN i67
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 43.605 26.885 44.175 ;
  END
 END i67
 PIN i68
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 39.425 26.885 39.995 ;
  END
 END i68
 PIN i69
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 35.435 26.885 36.005 ;
  END
 END i69
 PIN i70
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 31.255 26.885 31.825 ;
  END
 END i70
 PIN i71
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 689.415 26.885 689.985 ;
  END
 END i71
 PIN i72
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 27.265 26.885 27.835 ;
  END
 END i72
 PIN i73
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 23.085 26.885 23.655 ;
  END
 END i73
 PIN i74
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 19.095 26.885 19.665 ;
  END
 END i74
 PIN i75
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 14.915 26.885 15.485 ;
  END
 END i75
 PIN i76
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 10.925 26.885 11.495 ;
  END
 END i76
 PIN i77
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 6.745 26.885 7.315 ;
  END
 END i77
 PIN i78
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 2.755 26.885 3.325 ;
  END
 END i78
 PIN i79
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 685.425 26.885 685.995 ;
  END
 END i79
 PIN i80
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 681.245 26.885 681.815 ;
  END
 END i80
 PIN i81
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 677.255 26.885 677.825 ;
  END
 END i81
 PIN i82
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 673.075 26.885 673.645 ;
  END
 END i82
 PIN i83
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 742.615 26.885 743.185 ;
  END
 END i83
 PIN i84
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 650.845 26.885 651.415 ;
  END
 END i84
 PIN i85
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 646.665 26.885 647.235 ;
  END
 END i85
 PIN i86
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 642.675 26.885 643.245 ;
  END
 END i86
 PIN i87
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 638.495 26.885 639.065 ;
  END
 END i87
 PIN i88
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 634.505 26.885 635.075 ;
  END
 END i88
 PIN i89
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 630.325 26.885 630.895 ;
  END
 END i89
 PIN i90
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 626.335 26.885 626.905 ;
  END
 END i90
 PIN i91
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 622.155 26.885 622.725 ;
  END
 END i91
 PIN i92
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 618.165 26.885 618.735 ;
  END
 END i92
 PIN i93
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 613.985 26.885 614.555 ;
  END
 END i93
 PIN i94
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 738.435 26.885 739.005 ;
  END
 END i94
 PIN i95
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 609.995 26.885 610.565 ;
  END
 END i95
 PIN i96
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 605.815 26.885 606.385 ;
  END
 END i96
 PIN i97
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 601.825 26.885 602.395 ;
  END
 END i97
 PIN i98
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 597.645 26.885 598.215 ;
  END
 END i98
 PIN i99
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 593.655 26.885 594.225 ;
  END
 END i99
 PIN i100
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 589.475 26.885 590.045 ;
  END
 END i100
 PIN i101
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 585.485 26.885 586.055 ;
  END
 END i101
 PIN i102
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 581.305 26.885 581.875 ;
  END
 END i102
 PIN i103
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 577.315 26.885 577.885 ;
  END
 END i103
 PIN i104
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 573.135 26.885 573.705 ;
  END
 END i104
 PIN i105
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 734.445 26.885 735.015 ;
  END
 END i105
 PIN i106
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 564.015 26.885 564.585 ;
  END
 END i106
 PIN i107
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 559.835 26.885 560.405 ;
  END
 END i107
 PIN i108
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 555.845 26.885 556.415 ;
  END
 END i108
 PIN i109
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 551.665 26.885 552.235 ;
  END
 END i109
 PIN i110
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 547.675 26.885 548.245 ;
  END
 END i110
 PIN i111
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 543.495 26.885 544.065 ;
  END
 END i111
 PIN i112
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 539.505 26.885 540.075 ;
  END
 END i112
 PIN i113
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 535.325 26.885 535.895 ;
  END
 END i113
 PIN i114
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 531.335 26.885 531.905 ;
  END
 END i114
 PIN i115
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 527.155 26.885 527.725 ;
  END
 END i115
 PIN i116
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 730.265 26.885 730.835 ;
  END
 END i116
 PIN i117
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 523.165 26.885 523.735 ;
  END
 END i117
 PIN i118
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 518.985 26.885 519.555 ;
  END
 END i118
 PIN i119
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 514.995 26.885 515.565 ;
  END
 END i119
 PIN i120
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 510.815 26.885 511.385 ;
  END
 END i120
 PIN i121
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 506.825 26.885 507.395 ;
  END
 END i121
 PIN i122
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 502.645 26.885 503.215 ;
  END
 END i122
 PIN i123
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 498.655 26.885 499.225 ;
  END
 END i123
 PIN i124
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 494.475 26.885 495.045 ;
  END
 END i124
 PIN i125
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 490.485 26.885 491.055 ;
  END
 END i125
 PIN i126
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 486.305 26.885 486.875 ;
  END
 END i126
 PIN i127
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 726.275 26.885 726.845 ;
  END
 END i127
 PIN i128
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 464.075 26.885 464.645 ;
  END
 END i128
 PIN i129
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 459.895 26.885 460.465 ;
  END
 END i129
 PIN i130
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 455.905 26.885 456.475 ;
  END
 END i130
 PIN i131
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 451.725 26.885 452.295 ;
  END
 END i131
 PIN i132
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 447.735 26.885 448.305 ;
  END
 END i132
 PIN i133
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 443.555 26.885 444.125 ;
  END
 END i133
 PIN i134
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 439.565 26.885 440.135 ;
  END
 END i134
 PIN i135
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 435.385 26.885 435.955 ;
  END
 END i135
 PIN i136
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 431.395 26.885 431.965 ;
  END
 END i136
 PIN i137
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 427.215 26.885 427.785 ;
  END
 END i137
 PIN i138
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 722.095 26.885 722.665 ;
  END
 END i138
 PIN i139
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 423.225 26.885 423.795 ;
  END
 END i139
 PIN i140
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 419.045 26.885 419.615 ;
  END
 END i140
 PIN i141
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 415.055 26.885 415.625 ;
  END
 END i141
 PIN i142
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 410.875 26.885 411.445 ;
  END
 END i142
 PIN i143
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 406.885 26.885 407.455 ;
  END
 END i143
 PIN i144
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 402.705 26.885 403.275 ;
  END
 END i144
 PIN i145
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 398.715 26.885 399.285 ;
  END
 END i145
 PIN i146
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 394.535 26.885 395.105 ;
  END
 END i146
 PIN i147
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 390.545 26.885 391.115 ;
  END
 END i147
 PIN i148
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 386.365 26.885 386.935 ;
  END
 END i148
 PIN i149
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 718.105 26.885 718.675 ;
  END
 END i149
 PIN i150
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 354.825 26.885 355.395 ;
  END
 END i150
 PIN i151
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 350.645 26.885 351.215 ;
  END
 END i151
 PIN i152
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 346.655 26.885 347.225 ;
  END
 END i152
 PIN i153
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 342.475 26.885 343.045 ;
  END
 END i153
 PIN i154
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 338.485 26.885 339.055 ;
  END
 END i154
 PIN i155
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 334.305 26.885 334.875 ;
  END
 END i155
 PIN i156
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 330.315 26.885 330.885 ;
  END
 END i156
 PIN i157
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 326.135 26.885 326.705 ;
  END
 END i157
 PIN i158
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 322.145 26.885 322.715 ;
  END
 END i158
 PIN i159
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 317.965 26.885 318.535 ;
  END
 END i159
 PIN i160
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 713.925 26.885 714.495 ;
  END
 END i160
 PIN i161
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 313.975 26.885 314.545 ;
  END
 END i161
 PIN i162
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 309.795 26.885 310.365 ;
  END
 END i162
 PIN i163
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 305.805 26.885 306.375 ;
  END
 END i163
 PIN i164
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 301.625 26.885 302.195 ;
  END
 END i164
 PIN i165
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 297.635 26.885 298.205 ;
  END
 END i165
 PIN i166
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 293.455 26.885 294.025 ;
  END
 END i166
 PIN i167
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 289.465 26.885 290.035 ;
  END
 END i167
 PIN i168
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 285.285 26.885 285.855 ;
  END
 END i168
 PIN i169
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 281.295 26.885 281.865 ;
  END
 END i169
 PIN i170
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 277.115 26.885 277.685 ;
  END
 END i170
 PIN i171
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 695.305 27.645 695.875 ;
  END
 END i171
 PIN i172
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 691.315 27.645 691.885 ;
  END
 END i172
 PIN i173
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 687.135 27.645 687.705 ;
  END
 END i173
 PIN i174
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 707.655 27.645 708.225 ;
  END
 END i174
 PIN i175
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 703.475 27.645 704.045 ;
  END
 END i175
 PIN i176
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 628.045 27.645 628.615 ;
  END
 END i176
 PIN i177
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 624.055 27.645 624.625 ;
  END
 END i177
 PIN i178
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 619.875 27.645 620.445 ;
  END
 END i178
 PIN i179
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 615.885 27.645 616.455 ;
  END
 END i179
 PIN i180
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 611.705 27.645 612.275 ;
  END
 END i180
 PIN i181
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 508.535 27.645 509.105 ;
  END
 END i181
 PIN i182
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 504.545 27.645 505.115 ;
  END
 END i182
 PIN i183
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 500.365 27.645 500.935 ;
  END
 END i183
 PIN i184
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 520.885 27.645 521.455 ;
  END
 END i184
 PIN i185
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 516.705 27.645 517.275 ;
  END
 END i185
 PIN i186
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 441.275 27.645 441.845 ;
  END
 END i186
 PIN i187
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 437.285 27.645 437.855 ;
  END
 END i187
 PIN i188
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 433.105 27.645 433.675 ;
  END
 END i188
 PIN i189
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 429.115 27.645 429.685 ;
  END
 END i189
 PIN i190
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 424.935 27.645 425.505 ;
  END
 END i190
 PIN i191
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 299.915 27.645 300.485 ;
  END
 END i191
 PIN i192
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 303.905 27.645 304.475 ;
  END
 END i192
 PIN i193
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 308.085 27.645 308.655 ;
  END
 END i193
 PIN i194
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 312.075 27.645 312.645 ;
  END
 END i194
 PIN i195
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 316.255 27.645 316.825 ;
  END
 END i195
 PIN i196
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 232.655 27.645 233.225 ;
  END
 END i196
 PIN i197
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 236.645 27.645 237.215 ;
  END
 END i197
 PIN i198
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 240.825 27.645 241.395 ;
  END
 END i198
 PIN i199
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 220.305 27.645 220.875 ;
  END
 END i199
 PIN i200
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 224.485 27.645 225.055 ;
  END
 END i200
 PIN i201
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 121.315 27.645 121.885 ;
  END
 END i201
 PIN i202
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 125.305 27.645 125.875 ;
  END
 END i202
 PIN i203
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 129.485 27.645 130.055 ;
  END
 END i203
 PIN i204
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 133.475 27.645 134.045 ;
  END
 END i204
 PIN i205
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 137.655 27.645 138.225 ;
  END
 END i205
 PIN i206
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 54.055 27.645 54.625 ;
  END
 END i206
 PIN i207
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 58.045 27.645 58.615 ;
  END
 END i207
 PIN i208
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 62.225 27.645 62.795 ;
  END
 END i208
 PIN i209
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 41.705 27.645 42.275 ;
  END
 END i209
 PIN i210
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 45.885 27.645 46.455 ;
  END
 END i210
 PIN i211
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 699.485 27.645 700.055 ;
  END
 END i211
 PIN i212
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 632.225 27.645 632.795 ;
  END
 END i212
 PIN i213
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 512.715 27.645 513.285 ;
  END
 END i213
 PIN i214
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 445.455 27.645 446.025 ;
  END
 END i214
 PIN i215
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 295.735 27.645 296.305 ;
  END
 END i215
 PIN i216
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 228.475 27.645 229.045 ;
  END
 END i216
 PIN i217
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 117.135 27.645 117.705 ;
  END
 END i217
 PIN i218
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 49.875 27.645 50.445 ;
  END
 END i218
 PIN i219
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 17.955 382.945 18.525 383.515 ;
  END
 END i219
 PIN i220
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 17.955 369.645 18.525 370.215 ;
  END
 END i220
 PIN i221
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 750.215 27.645 750.785 ;
  END
 END i221
 PIN i222
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 746.035 27.645 746.605 ;
  END
 END i222
 PIN i223
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 709.365 27.645 709.935 ;
  END
 END i223
 PIN i224
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 255.455 27.645 256.025 ;
  END
 END i224
 PIN i225
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 251.275 27.645 251.845 ;
  END
 END i225
 PIN i226
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 247.285 27.645 247.855 ;
  END
 END i226
 PIN i227
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 243.105 27.645 243.675 ;
  END
 END i227
 PIN i228
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 239.115 27.645 239.685 ;
  END
 END i228
 PIN i229
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 234.935 27.645 235.505 ;
  END
 END i229
 PIN i230
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 230.945 27.645 231.515 ;
  END
 END i230
 PIN i231
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 226.765 27.645 227.335 ;
  END
 END i231
 PIN i232
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 222.775 27.645 223.345 ;
  END
 END i232
 PIN i233
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 218.595 27.645 219.165 ;
  END
 END i233
 PIN i234
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 705.185 27.645 705.755 ;
  END
 END i234
 PIN i235
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 214.605 27.645 215.175 ;
  END
 END i235
 PIN i236
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 210.425 27.645 210.995 ;
  END
 END i236
 PIN i237
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 206.435 27.645 207.005 ;
  END
 END i237
 PIN i238
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 202.255 27.645 202.825 ;
  END
 END i238
 PIN i239
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 198.265 27.645 198.835 ;
  END
 END i239
 PIN i240
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 194.085 27.645 194.655 ;
  END
 END i240
 PIN i241
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 190.095 27.645 190.665 ;
  END
 END i241
 PIN i242
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 185.915 27.645 186.485 ;
  END
 END i242
 PIN i243
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 181.925 27.645 182.495 ;
  END
 END i243
 PIN i244
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 172.615 27.645 173.185 ;
  END
 END i244
 PIN i245
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 701.195 27.645 701.765 ;
  END
 END i245
 PIN i246
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 168.625 27.645 169.195 ;
  END
 END i246
 PIN i247
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 164.445 27.645 165.015 ;
  END
 END i247
 PIN i248
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 160.455 27.645 161.025 ;
  END
 END i248
 PIN i249
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 156.275 27.645 156.845 ;
  END
 END i249
 PIN i250
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 152.285 27.645 152.855 ;
  END
 END i250
 PIN i251
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 148.105 27.645 148.675 ;
  END
 END i251
 PIN i252
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 144.115 27.645 144.685 ;
  END
 END i252
 PIN i253
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 139.935 27.645 140.505 ;
  END
 END i253
 PIN i254
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 135.945 27.645 136.515 ;
  END
 END i254
 PIN i255
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 131.765 27.645 132.335 ;
  END
 END i255
 PIN i256
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 697.015 27.645 697.585 ;
  END
 END i256
 PIN i257
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 127.775 27.645 128.345 ;
  END
 END i257
 PIN i258
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 123.595 27.645 124.165 ;
  END
 END i258
 PIN i259
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 119.605 27.645 120.175 ;
  END
 END i259
 PIN i260
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 115.425 27.645 115.995 ;
  END
 END i260
 PIN i261
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 111.435 27.645 112.005 ;
  END
 END i261
 PIN i262
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 107.255 27.645 107.825 ;
  END
 END i262
 PIN i263
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 103.265 27.645 103.835 ;
  END
 END i263
 PIN i264
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 99.085 27.645 99.655 ;
  END
 END i264
 PIN i265
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 76.855 27.645 77.425 ;
  END
 END i265
 PIN i266
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 72.675 27.645 73.245 ;
  END
 END i266
 PIN i267
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 693.025 27.645 693.595 ;
  END
 END i267
 PIN i268
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 68.685 27.645 69.255 ;
  END
 END i268
 PIN i269
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 64.505 27.645 65.075 ;
  END
 END i269
 PIN i270
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 60.515 27.645 61.085 ;
  END
 END i270
 PIN i271
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 56.335 27.645 56.905 ;
  END
 END i271
 PIN i272
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 52.345 27.645 52.915 ;
  END
 END i272
 PIN i273
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 48.165 27.645 48.735 ;
  END
 END i273
 PIN i274
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 44.175 27.645 44.745 ;
  END
 END i274
 PIN i275
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 39.995 27.645 40.565 ;
  END
 END i275
 PIN i276
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 36.005 27.645 36.575 ;
  END
 END i276
 PIN i277
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 31.825 27.645 32.395 ;
  END
 END i277
 PIN i278
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 688.845 27.645 689.415 ;
  END
 END i278
 PIN i279
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 27.835 27.645 28.405 ;
  END
 END i279
 PIN i280
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 23.655 27.645 24.225 ;
  END
 END i280
 PIN i281
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 19.665 27.645 20.235 ;
  END
 END i281
 PIN i282
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 15.485 27.645 16.055 ;
  END
 END i282
 PIN i283
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 11.495 27.645 12.065 ;
  END
 END i283
 PIN i284
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 7.315 27.645 7.885 ;
  END
 END i284
 PIN i285
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 3.325 27.645 3.895 ;
  END
 END i285
 PIN i286
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 684.855 27.645 685.425 ;
  END
 END i286
 PIN i287
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 680.675 27.645 681.245 ;
  END
 END i287
 PIN i288
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 676.685 27.645 677.255 ;
  END
 END i288
 PIN i289
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 672.505 27.645 673.075 ;
  END
 END i289
 PIN i290
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 742.045 27.645 742.615 ;
  END
 END i290
 PIN i291
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 650.275 27.645 650.845 ;
  END
 END i291
 PIN i292
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 646.095 27.645 646.665 ;
  END
 END i292
 PIN i293
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 642.105 27.645 642.675 ;
  END
 END i293
 PIN i294
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 637.925 27.645 638.495 ;
  END
 END i294
 PIN i295
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 633.935 27.645 634.505 ;
  END
 END i295
 PIN i296
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 629.755 27.645 630.325 ;
  END
 END i296
 PIN i297
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 625.765 27.645 626.335 ;
  END
 END i297
 PIN i298
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 621.585 27.645 622.155 ;
  END
 END i298
 PIN i299
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 617.595 27.645 618.165 ;
  END
 END i299
 PIN i300
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 613.415 27.645 613.985 ;
  END
 END i300
 PIN i301
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 737.865 27.645 738.435 ;
  END
 END i301
 PIN i302
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 609.425 27.645 609.995 ;
  END
 END i302
 PIN i303
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 605.245 27.645 605.815 ;
  END
 END i303
 PIN i304
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 601.255 27.645 601.825 ;
  END
 END i304
 PIN i305
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 597.075 27.645 597.645 ;
  END
 END i305
 PIN i306
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 593.085 27.645 593.655 ;
  END
 END i306
 PIN i307
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 588.905 27.645 589.475 ;
  END
 END i307
 PIN i308
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 584.915 27.645 585.485 ;
  END
 END i308
 PIN i309
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 580.735 27.645 581.305 ;
  END
 END i309
 PIN i310
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 576.745 27.645 577.315 ;
  END
 END i310
 PIN i311
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 572.565 27.645 573.135 ;
  END
 END i311
 PIN i312
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 733.875 27.645 734.445 ;
  END
 END i312
 PIN i313
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 563.445 27.645 564.015 ;
  END
 END i313
 PIN i314
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 559.265 27.645 559.835 ;
  END
 END i314
 PIN i315
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 555.275 27.645 555.845 ;
  END
 END i315
 PIN i316
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 551.095 27.645 551.665 ;
  END
 END i316
 PIN i317
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 547.105 27.645 547.675 ;
  END
 END i317
 PIN i318
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 542.925 27.645 543.495 ;
  END
 END i318
 PIN i319
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 538.935 27.645 539.505 ;
  END
 END i319
 PIN i320
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 534.755 27.645 535.325 ;
  END
 END i320
 PIN i321
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 530.765 27.645 531.335 ;
  END
 END i321
 PIN i322
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 526.585 27.645 527.155 ;
  END
 END i322
 PIN i323
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 729.695 27.645 730.265 ;
  END
 END i323
 PIN i324
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 522.595 27.645 523.165 ;
  END
 END i324
 PIN i325
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 518.415 27.645 518.985 ;
  END
 END i325
 PIN i326
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 514.425 27.645 514.995 ;
  END
 END i326
 PIN i327
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 510.245 27.645 510.815 ;
  END
 END i327
 PIN i328
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 506.255 27.645 506.825 ;
  END
 END i328
 PIN i329
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 502.075 27.645 502.645 ;
  END
 END i329
 PIN i330
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 498.085 27.645 498.655 ;
  END
 END i330
 PIN i331
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 493.905 27.645 494.475 ;
  END
 END i331
 PIN i332
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 489.915 27.645 490.485 ;
  END
 END i332
 PIN i333
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 485.735 27.645 486.305 ;
  END
 END i333
 PIN i334
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 725.705 27.645 726.275 ;
  END
 END i334
 PIN i335
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 463.505 27.645 464.075 ;
  END
 END i335
 PIN i336
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 459.325 27.645 459.895 ;
  END
 END i336
 PIN i337
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 455.335 27.645 455.905 ;
  END
 END i337
 PIN i338
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 451.155 27.645 451.725 ;
  END
 END i338
 PIN i339
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 447.165 27.645 447.735 ;
  END
 END i339
 PIN i340
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 442.985 27.645 443.555 ;
  END
 END i340
 PIN i341
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 438.995 27.645 439.565 ;
  END
 END i341
 PIN i342
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 434.815 27.645 435.385 ;
  END
 END i342
 PIN i343
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 430.825 27.645 431.395 ;
  END
 END i343
 PIN i344
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 426.645 27.645 427.215 ;
  END
 END i344
 PIN i345
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 721.525 27.645 722.095 ;
  END
 END i345
 PIN i346
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 422.655 27.645 423.225 ;
  END
 END i346
 PIN i347
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 418.475 27.645 419.045 ;
  END
 END i347
 PIN i348
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 414.485 27.645 415.055 ;
  END
 END i348
 PIN i349
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 410.305 27.645 410.875 ;
  END
 END i349
 PIN i350
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 406.315 27.645 406.885 ;
  END
 END i350
 PIN i351
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 402.135 27.645 402.705 ;
  END
 END i351
 PIN i352
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 398.145 27.645 398.715 ;
  END
 END i352
 PIN i353
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 393.965 27.645 394.535 ;
  END
 END i353
 PIN i354
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 389.975 27.645 390.545 ;
  END
 END i354
 PIN i355
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 385.795 27.645 386.365 ;
  END
 END i355
 PIN i356
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 717.535 27.645 718.105 ;
  END
 END i356
 PIN i357
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 355.395 27.645 355.965 ;
  END
 END i357
 PIN i358
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 351.215 27.645 351.785 ;
  END
 END i358
 PIN i359
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 347.225 27.645 347.795 ;
  END
 END i359
 PIN i360
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 343.045 27.645 343.615 ;
  END
 END i360
 PIN i361
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 339.055 27.645 339.625 ;
  END
 END i361
 PIN i362
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 334.875 27.645 335.445 ;
  END
 END i362
 PIN i363
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 330.885 27.645 331.455 ;
  END
 END i363
 PIN i364
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 326.705 27.645 327.275 ;
  END
 END i364
 PIN i365
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 322.715 27.645 323.285 ;
  END
 END i365
 PIN i366
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 318.535 27.645 319.105 ;
  END
 END i366
 PIN i367
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 713.355 27.645 713.925 ;
  END
 END i367
 PIN i368
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 314.545 27.645 315.115 ;
  END
 END i368
 PIN i369
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 310.365 27.645 310.935 ;
  END
 END i369
 PIN i370
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 306.375 27.645 306.945 ;
  END
 END i370
 PIN i371
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 302.195 27.645 302.765 ;
  END
 END i371
 PIN i372
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 298.205 27.645 298.775 ;
  END
 END i372
 PIN i373
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 294.025 27.645 294.595 ;
  END
 END i373
 PIN i374
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 290.035 27.645 290.605 ;
  END
 END i374
 PIN i375
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 285.855 27.645 286.425 ;
  END
 END i375
 PIN i376
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 281.865 27.645 282.435 ;
  END
 END i376
 PIN i377
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 277.685 27.645 278.255 ;
  END
 END i377
 PIN i378
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 375.345 3.705 375.915 ;
  END
 END i378
 PIN i379
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 374.965 4.465 375.535 ;
  END
 END i379
 PIN i380
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 749.645 28.405 750.215 ;
  END
 END i380
 PIN i381
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 745.465 28.405 746.035 ;
  END
 END i381
 PIN i382
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 708.795 28.405 709.365 ;
  END
 END i382
 PIN i383
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 256.025 28.405 256.595 ;
  END
 END i383
 PIN i384
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 251.845 28.405 252.415 ;
  END
 END i384
 PIN i385
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 247.855 28.405 248.425 ;
  END
 END i385
 PIN i386
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 243.675 28.405 244.245 ;
  END
 END i386
 PIN i387
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 239.685 28.405 240.255 ;
  END
 END i387
 PIN i388
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 235.505 28.405 236.075 ;
  END
 END i388
 PIN i389
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 231.515 28.405 232.085 ;
  END
 END i389
 PIN i390
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 227.335 28.405 227.905 ;
  END
 END i390
 PIN i391
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 223.345 28.405 223.915 ;
  END
 END i391
 PIN i392
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 219.165 28.405 219.735 ;
  END
 END i392
 PIN i393
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 704.615 28.405 705.185 ;
  END
 END i393
 PIN i394
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 215.175 28.405 215.745 ;
  END
 END i394
 PIN i395
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 210.995 28.405 211.565 ;
  END
 END i395
 PIN i396
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 207.005 28.405 207.575 ;
  END
 END i396
 PIN i397
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 202.825 28.405 203.395 ;
  END
 END i397
 PIN i398
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 198.835 28.405 199.405 ;
  END
 END i398
 PIN i399
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 194.655 28.405 195.225 ;
  END
 END i399
 PIN i400
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 190.665 28.405 191.235 ;
  END
 END i400
 PIN i401
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 186.485 28.405 187.055 ;
  END
 END i401
 PIN i402
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 182.495 28.405 183.065 ;
  END
 END i402
 PIN i403
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 173.185 28.405 173.755 ;
  END
 END i403
 PIN i404
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 700.625 28.405 701.195 ;
  END
 END i404
 PIN i405
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 169.195 28.405 169.765 ;
  END
 END i405
 PIN i406
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 165.015 28.405 165.585 ;
  END
 END i406
 PIN i407
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 161.025 28.405 161.595 ;
  END
 END i407
 PIN i408
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 156.845 28.405 157.415 ;
  END
 END i408
 PIN i409
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 152.855 28.405 153.425 ;
  END
 END i409
 PIN i410
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 148.675 28.405 149.245 ;
  END
 END i410
 PIN i411
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 144.685 28.405 145.255 ;
  END
 END i411
 PIN i412
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 140.505 28.405 141.075 ;
  END
 END i412
 PIN i413
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 136.515 28.405 137.085 ;
  END
 END i413
 PIN i414
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 132.335 28.405 132.905 ;
  END
 END i414
 PIN i415
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 696.445 28.405 697.015 ;
  END
 END i415
 PIN i416
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 128.345 28.405 128.915 ;
  END
 END i416
 PIN i417
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 124.165 28.405 124.735 ;
  END
 END i417
 PIN i418
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 120.175 28.405 120.745 ;
  END
 END i418
 PIN i419
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 115.995 28.405 116.565 ;
  END
 END i419
 PIN i420
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 112.005 28.405 112.575 ;
  END
 END i420
 PIN i421
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 107.825 28.405 108.395 ;
  END
 END i421
 PIN i422
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 103.835 28.405 104.405 ;
  END
 END i422
 PIN i423
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 99.655 28.405 100.225 ;
  END
 END i423
 PIN i424
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 77.425 28.405 77.995 ;
  END
 END i424
 PIN i425
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 73.245 28.405 73.815 ;
  END
 END i425
 PIN i426
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 692.455 28.405 693.025 ;
  END
 END i426
 PIN i427
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 69.255 28.405 69.825 ;
  END
 END i427
 PIN i428
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 65.075 28.405 65.645 ;
  END
 END i428
 PIN i429
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 61.085 28.405 61.655 ;
  END
 END i429
 PIN i430
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 56.905 28.405 57.475 ;
  END
 END i430
 PIN i431
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 52.915 28.405 53.485 ;
  END
 END i431
 PIN i432
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 48.735 28.405 49.305 ;
  END
 END i432
 PIN i433
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 44.745 28.405 45.315 ;
  END
 END i433
 PIN i434
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 40.565 28.405 41.135 ;
  END
 END i434
 PIN i435
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 36.575 28.405 37.145 ;
  END
 END i435
 PIN i436
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 32.395 28.405 32.965 ;
  END
 END i436
 PIN i437
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 688.275 28.405 688.845 ;
  END
 END i437
 PIN i438
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 28.405 28.405 28.975 ;
  END
 END i438
 PIN i439
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 24.225 28.405 24.795 ;
  END
 END i439
 PIN i440
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 20.235 28.405 20.805 ;
  END
 END i440
 PIN i441
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 16.055 28.405 16.625 ;
  END
 END i441
 PIN i442
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 12.065 28.405 12.635 ;
  END
 END i442
 PIN i443
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 7.885 28.405 8.455 ;
  END
 END i443
 PIN i444
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 3.895 28.405 4.465 ;
  END
 END i444
 PIN i445
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 684.285 28.405 684.855 ;
  END
 END i445
 PIN i446
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 680.105 28.405 680.675 ;
  END
 END i446
 PIN i447
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 676.115 28.405 676.685 ;
  END
 END i447
 PIN i448
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 671.935 28.405 672.505 ;
  END
 END i448
 PIN i449
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 741.475 28.405 742.045 ;
  END
 END i449
 PIN i450
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 649.705 28.405 650.275 ;
  END
 END i450
 PIN i451
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 645.525 28.405 646.095 ;
  END
 END i451
 PIN i452
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 641.535 28.405 642.105 ;
  END
 END i452
 PIN i453
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 637.355 28.405 637.925 ;
  END
 END i453
 PIN i454
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 633.365 28.405 633.935 ;
  END
 END i454
 PIN i455
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 629.185 28.405 629.755 ;
  END
 END i455
 PIN i456
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 625.195 28.405 625.765 ;
  END
 END i456
 PIN i457
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 621.015 28.405 621.585 ;
  END
 END i457
 PIN i458
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 617.025 28.405 617.595 ;
  END
 END i458
 PIN i459
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 612.845 28.405 613.415 ;
  END
 END i459
 PIN i460
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 737.295 28.405 737.865 ;
  END
 END i460
 PIN i461
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 608.855 28.405 609.425 ;
  END
 END i461
 PIN i462
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 604.675 28.405 605.245 ;
  END
 END i462
 PIN i463
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 600.685 28.405 601.255 ;
  END
 END i463
 PIN i464
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 596.505 28.405 597.075 ;
  END
 END i464
 PIN i465
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 592.515 28.405 593.085 ;
  END
 END i465
 PIN i466
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 588.335 28.405 588.905 ;
  END
 END i466
 PIN i467
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 584.345 28.405 584.915 ;
  END
 END i467
 PIN i468
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 580.165 28.405 580.735 ;
  END
 END i468
 PIN i469
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 576.175 28.405 576.745 ;
  END
 END i469
 PIN i470
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 571.995 28.405 572.565 ;
  END
 END i470
 PIN i471
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 733.305 28.405 733.875 ;
  END
 END i471
 PIN i472
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 562.875 28.405 563.445 ;
  END
 END i472
 PIN i473
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 558.695 28.405 559.265 ;
  END
 END i473
 PIN i474
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 554.705 28.405 555.275 ;
  END
 END i474
 PIN i475
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 550.525 28.405 551.095 ;
  END
 END i475
 PIN i476
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 546.535 28.405 547.105 ;
  END
 END i476
 PIN i477
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 542.355 28.405 542.925 ;
  END
 END i477
 PIN i478
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 538.365 28.405 538.935 ;
  END
 END i478
 PIN i479
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 534.185 28.405 534.755 ;
  END
 END i479
 PIN i480
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 530.195 28.405 530.765 ;
  END
 END i480
 PIN i481
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 526.015 28.405 526.585 ;
  END
 END i481
 PIN i482
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 729.125 28.405 729.695 ;
  END
 END i482
 PIN i483
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 522.025 28.405 522.595 ;
  END
 END i483
 PIN i484
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 517.845 28.405 518.415 ;
  END
 END i484
 PIN i485
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 513.855 28.405 514.425 ;
  END
 END i485
 PIN i486
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 509.675 28.405 510.245 ;
  END
 END i486
 PIN i487
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 505.685 28.405 506.255 ;
  END
 END i487
 PIN i488
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 501.505 28.405 502.075 ;
  END
 END i488
 PIN i489
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 497.515 28.405 498.085 ;
  END
 END i489
 PIN i490
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 493.335 28.405 493.905 ;
  END
 END i490
 PIN i491
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 489.345 28.405 489.915 ;
  END
 END i491
 PIN i492
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 485.165 28.405 485.735 ;
  END
 END i492
 PIN i493
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 725.135 28.405 725.705 ;
  END
 END i493
 PIN i494
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 462.935 28.405 463.505 ;
  END
 END i494
 PIN i495
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 458.755 28.405 459.325 ;
  END
 END i495
 PIN i496
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 454.765 28.405 455.335 ;
  END
 END i496
 PIN i497
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 450.585 28.405 451.155 ;
  END
 END i497
 PIN i498
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 446.595 28.405 447.165 ;
  END
 END i498
 PIN i499
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 442.415 28.405 442.985 ;
  END
 END i499
 PIN i500
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 438.425 28.405 438.995 ;
  END
 END i500
 PIN i501
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 434.245 28.405 434.815 ;
  END
 END i501
 PIN i502
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 430.255 28.405 430.825 ;
  END
 END i502
 PIN i503
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 426.075 28.405 426.645 ;
  END
 END i503
 PIN i504
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 720.955 28.405 721.525 ;
  END
 END i504
 PIN i505
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 422.085 28.405 422.655 ;
  END
 END i505
 PIN i506
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 417.905 28.405 418.475 ;
  END
 END i506
 PIN i507
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 413.915 28.405 414.485 ;
  END
 END i507
 PIN i508
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 409.735 28.405 410.305 ;
  END
 END i508
 PIN i509
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 405.745 28.405 406.315 ;
  END
 END i509
 PIN i510
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 401.565 28.405 402.135 ;
  END
 END i510
 PIN i511
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 397.575 28.405 398.145 ;
  END
 END i511
 PIN i512
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 393.395 28.405 393.965 ;
  END
 END i512
 PIN i513
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 389.405 28.405 389.975 ;
  END
 END i513
 PIN i514
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 385.225 28.405 385.795 ;
  END
 END i514
 PIN i515
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 716.965 28.405 717.535 ;
  END
 END i515
 PIN i516
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 355.965 28.405 356.535 ;
  END
 END i516
 PIN i517
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 351.785 28.405 352.355 ;
  END
 END i517
 PIN i518
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 347.795 28.405 348.365 ;
  END
 END i518
 PIN i519
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 343.615 28.405 344.185 ;
  END
 END i519
 PIN i520
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 339.625 28.405 340.195 ;
  END
 END i520
 PIN i521
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 335.445 28.405 336.015 ;
  END
 END i521
 PIN i522
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 331.455 28.405 332.025 ;
  END
 END i522
 PIN i523
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 327.275 28.405 327.845 ;
  END
 END i523
 PIN i524
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 323.285 28.405 323.855 ;
  END
 END i524
 PIN i525
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 319.105 28.405 319.675 ;
  END
 END i525
 PIN i526
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 712.785 28.405 713.355 ;
  END
 END i526
 PIN i527
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 315.115 28.405 315.685 ;
  END
 END i527
 PIN i528
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 310.935 28.405 311.505 ;
  END
 END i528
 PIN i529
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 306.945 28.405 307.515 ;
  END
 END i529
 PIN i530
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 302.765 28.405 303.335 ;
  END
 END i530
 PIN i531
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 298.775 28.405 299.345 ;
  END
 END i531
 PIN i532
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 294.595 28.405 295.165 ;
  END
 END i532
 PIN i533
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 290.605 28.405 291.175 ;
  END
 END i533
 PIN i534
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 286.425 28.405 286.995 ;
  END
 END i534
 PIN i535
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 282.435 28.405 283.005 ;
  END
 END i535
 PIN i536
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 278.255 28.405 278.825 ;
  END
 END i536
 PIN i537
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 4.275 382.945 4.845 383.515 ;
  END
 END i537
 PIN i538
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 5.415 382.945 5.985 383.515 ;
  END
 END i538
 PIN i539
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 6.935 382.945 7.505 383.515 ;
  END
 END i539
 PIN i540
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 8.835 382.945 9.405 383.515 ;
  END
 END i540
 PIN i541
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 4.275 369.645 4.845 370.215 ;
  END
 END i541
 PIN i542
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 5.415 369.645 5.985 370.215 ;
  END
 END i542
 PIN i543
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 6.935 369.645 7.505 370.215 ;
  END
 END i543
 PIN i544
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 8.835 369.645 9.405 370.215 ;
  END
 END i544
 OBS
  LAYER metal1 ;
   RECT 23.18 0.0 157.32 1.71 ;
   RECT 23.18 1.71 157.32 3.42 ;
   RECT 23.18 3.42 157.32 5.13 ;
   RECT 23.18 5.13 157.32 6.84 ;
   RECT 23.18 6.84 157.32 8.55 ;
   RECT 23.18 8.55 157.32 10.26 ;
   RECT 23.18 10.26 157.32 11.97 ;
   RECT 23.18 11.97 157.32 13.68 ;
   RECT 23.18 13.68 157.32 15.39 ;
   RECT 23.18 15.39 157.32 17.1 ;
   RECT 23.18 17.1 157.32 18.81 ;
   RECT 23.18 18.81 157.32 20.52 ;
   RECT 23.18 20.52 157.32 22.23 ;
   RECT 23.18 22.23 157.32 23.94 ;
   RECT 23.18 23.94 157.32 25.65 ;
   RECT 23.18 25.65 157.32 27.36 ;
   RECT 23.18 27.36 157.32 29.07 ;
   RECT 23.18 29.07 157.32 30.78 ;
   RECT 23.18 30.78 157.32 32.49 ;
   RECT 23.18 32.49 157.32 34.2 ;
   RECT 23.18 34.2 157.32 35.91 ;
   RECT 23.18 35.91 157.32 37.62 ;
   RECT 23.18 37.62 157.32 39.33 ;
   RECT 23.18 39.33 157.32 41.04 ;
   RECT 23.18 41.04 157.32 42.75 ;
   RECT 23.18 42.75 157.32 44.46 ;
   RECT 23.18 44.46 157.32 46.17 ;
   RECT 23.18 46.17 157.32 47.88 ;
   RECT 23.18 47.88 157.32 49.59 ;
   RECT 23.18 49.59 157.32 51.3 ;
   RECT 23.18 51.3 157.32 53.01 ;
   RECT 23.18 53.01 157.32 54.72 ;
   RECT 23.18 54.72 157.32 56.43 ;
   RECT 23.18 56.43 157.32 58.14 ;
   RECT 23.18 58.14 157.32 59.85 ;
   RECT 23.18 59.85 157.32 61.56 ;
   RECT 23.18 61.56 157.32 63.27 ;
   RECT 23.18 63.27 157.32 64.98 ;
   RECT 23.18 64.98 157.32 66.69 ;
   RECT 23.18 66.69 157.32 68.4 ;
   RECT 23.18 68.4 157.32 70.11 ;
   RECT 23.18 70.11 157.32 71.82 ;
   RECT 23.18 71.82 157.32 73.53 ;
   RECT 23.18 73.53 157.32 75.24 ;
   RECT 23.18 75.24 157.32 76.95 ;
   RECT 23.18 76.95 157.32 78.66 ;
   RECT 23.18 78.66 157.32 80.37 ;
   RECT 23.18 80.37 157.32 82.08 ;
   RECT 23.18 82.08 157.32 83.79 ;
   RECT 23.18 83.79 157.32 85.5 ;
   RECT 23.18 85.5 157.32 87.21 ;
   RECT 23.18 87.21 157.32 88.92 ;
   RECT 23.18 88.92 157.32 90.63 ;
   RECT 23.18 90.63 157.32 92.34 ;
   RECT 23.18 92.34 157.32 94.05 ;
   RECT 23.18 94.05 157.32 95.76 ;
   RECT 23.18 95.76 157.32 97.47 ;
   RECT 23.18 97.47 157.32 99.18 ;
   RECT 23.18 99.18 157.32 100.89 ;
   RECT 23.18 100.89 157.32 102.6 ;
   RECT 23.18 102.6 157.32 104.31 ;
   RECT 23.18 104.31 157.32 106.02 ;
   RECT 23.18 106.02 157.32 107.73 ;
   RECT 23.18 107.73 157.32 109.44 ;
   RECT 23.18 109.44 157.32 111.15 ;
   RECT 23.18 111.15 157.32 112.86 ;
   RECT 23.18 112.86 157.32 114.57 ;
   RECT 23.18 114.57 157.32 116.28 ;
   RECT 23.18 116.28 157.32 117.99 ;
   RECT 23.18 117.99 157.32 119.7 ;
   RECT 23.18 119.7 157.32 121.41 ;
   RECT 23.18 121.41 157.32 123.12 ;
   RECT 23.18 123.12 157.32 124.83 ;
   RECT 23.18 124.83 157.32 126.54 ;
   RECT 23.18 126.54 157.32 128.25 ;
   RECT 23.18 128.25 157.32 129.96 ;
   RECT 23.18 129.96 157.32 131.67 ;
   RECT 23.18 131.67 157.32 133.38 ;
   RECT 23.18 133.38 157.32 135.09 ;
   RECT 23.18 135.09 157.32 136.8 ;
   RECT 23.18 136.8 157.32 138.51 ;
   RECT 23.18 138.51 157.32 140.22 ;
   RECT 23.18 140.22 157.32 141.93 ;
   RECT 23.18 141.93 157.32 143.64 ;
   RECT 23.18 143.64 157.32 145.35 ;
   RECT 23.18 145.35 157.32 147.06 ;
   RECT 23.18 147.06 157.32 148.77 ;
   RECT 23.18 148.77 157.32 150.48 ;
   RECT 23.18 150.48 157.32 152.19 ;
   RECT 23.18 152.19 157.32 153.9 ;
   RECT 23.18 153.9 157.32 155.61 ;
   RECT 23.18 155.61 157.32 157.32 ;
   RECT 23.18 157.32 157.32 159.03 ;
   RECT 23.18 159.03 157.32 160.74 ;
   RECT 23.18 160.74 157.32 162.45 ;
   RECT 23.18 162.45 157.32 164.16 ;
   RECT 23.18 164.16 157.32 165.87 ;
   RECT 23.18 165.87 157.32 167.58 ;
   RECT 23.18 167.58 157.32 169.29 ;
   RECT 23.18 169.29 157.32 171.0 ;
   RECT 23.18 171.0 157.32 172.71 ;
   RECT 23.18 172.71 157.32 174.42 ;
   RECT 23.18 174.42 157.32 176.13 ;
   RECT 23.18 176.13 157.32 177.84 ;
   RECT 23.18 177.84 157.32 179.55 ;
   RECT 23.18 179.55 157.32 181.26 ;
   RECT 23.18 181.26 157.32 182.97 ;
   RECT 23.18 182.97 157.32 184.68 ;
   RECT 23.18 184.68 157.32 186.39 ;
   RECT 23.18 186.39 157.32 188.1 ;
   RECT 23.18 188.1 157.32 189.81 ;
   RECT 23.18 189.81 157.32 191.52 ;
   RECT 23.18 191.52 157.32 193.23 ;
   RECT 23.18 193.23 157.32 194.94 ;
   RECT 23.18 194.94 157.32 196.65 ;
   RECT 23.18 196.65 157.32 198.36 ;
   RECT 23.18 198.36 157.32 200.07 ;
   RECT 23.18 200.07 157.32 201.78 ;
   RECT 23.18 201.78 157.32 203.49 ;
   RECT 23.18 203.49 157.32 205.2 ;
   RECT 23.18 205.2 157.32 206.91 ;
   RECT 23.18 206.91 157.32 208.62 ;
   RECT 23.18 208.62 157.32 210.33 ;
   RECT 23.18 210.33 157.32 212.04 ;
   RECT 23.18 212.04 157.32 213.75 ;
   RECT 23.18 213.75 157.32 215.46 ;
   RECT 23.18 215.46 157.32 217.17 ;
   RECT 23.18 217.17 157.32 218.88 ;
   RECT 23.18 218.88 157.32 220.59 ;
   RECT 23.18 220.59 157.32 222.3 ;
   RECT 23.18 222.3 157.32 224.01 ;
   RECT 23.18 224.01 157.32 225.72 ;
   RECT 23.18 225.72 157.32 227.43 ;
   RECT 23.18 227.43 157.32 229.14 ;
   RECT 23.18 229.14 157.32 230.85 ;
   RECT 23.18 230.85 157.32 232.56 ;
   RECT 23.18 232.56 157.32 234.27 ;
   RECT 23.18 234.27 157.32 235.98 ;
   RECT 23.18 235.98 157.32 237.69 ;
   RECT 23.18 237.69 157.32 239.4 ;
   RECT 23.18 239.4 157.32 241.11 ;
   RECT 23.18 241.11 157.32 242.82 ;
   RECT 23.18 242.82 157.32 244.53 ;
   RECT 23.18 244.53 157.32 246.24 ;
   RECT 23.18 246.24 157.32 247.95 ;
   RECT 23.18 247.95 157.32 249.66 ;
   RECT 23.18 249.66 157.32 251.37 ;
   RECT 23.18 251.37 157.32 253.08 ;
   RECT 23.18 253.08 157.32 254.79 ;
   RECT 23.18 254.79 157.32 256.5 ;
   RECT 23.18 256.5 157.32 258.21 ;
   RECT 23.18 258.21 157.32 259.92 ;
   RECT 23.18 259.92 157.32 261.63 ;
   RECT 23.18 261.63 157.32 263.34 ;
   RECT 23.18 263.34 157.32 265.05 ;
   RECT 23.18 265.05 157.32 266.76 ;
   RECT 23.18 266.76 157.32 268.47 ;
   RECT 23.18 268.47 157.32 270.18 ;
   RECT 23.18 270.18 157.32 271.89 ;
   RECT 23.18 271.89 157.32 273.6 ;
   RECT 23.18 273.6 157.32 275.31 ;
   RECT 23.18 275.31 157.32 277.02 ;
   RECT 23.18 277.02 157.32 278.73 ;
   RECT 23.18 278.73 157.32 280.44 ;
   RECT 23.18 280.44 157.32 282.15 ;
   RECT 23.18 282.15 157.32 283.86 ;
   RECT 23.18 283.86 157.32 285.57 ;
   RECT 23.18 285.57 157.32 287.28 ;
   RECT 23.18 287.28 157.32 288.99 ;
   RECT 23.18 288.99 157.32 290.7 ;
   RECT 23.18 290.7 157.32 292.41 ;
   RECT 23.18 292.41 157.32 294.12 ;
   RECT 23.18 294.12 157.32 295.83 ;
   RECT 23.18 295.83 157.32 297.54 ;
   RECT 23.18 297.54 157.32 299.25 ;
   RECT 23.18 299.25 157.32 300.96 ;
   RECT 23.18 300.96 157.32 302.67 ;
   RECT 23.18 302.67 157.32 304.38 ;
   RECT 23.18 304.38 157.32 306.09 ;
   RECT 23.18 306.09 157.32 307.8 ;
   RECT 23.18 307.8 157.32 309.51 ;
   RECT 23.18 309.51 157.32 311.22 ;
   RECT 23.18 311.22 157.32 312.93 ;
   RECT 23.18 312.93 157.32 314.64 ;
   RECT 23.18 314.64 157.32 316.35 ;
   RECT 23.18 316.35 157.32 318.06 ;
   RECT 23.18 318.06 157.32 319.77 ;
   RECT 23.18 319.77 157.32 321.48 ;
   RECT 23.18 321.48 157.32 323.19 ;
   RECT 23.18 323.19 157.32 324.9 ;
   RECT 23.18 324.9 157.32 326.61 ;
   RECT 23.18 326.61 157.32 328.32 ;
   RECT 23.18 328.32 157.32 330.03 ;
   RECT 23.18 330.03 157.32 331.74 ;
   RECT 23.18 331.74 157.32 333.45 ;
   RECT 23.18 333.45 157.32 335.16 ;
   RECT 23.18 335.16 157.32 336.87 ;
   RECT 23.18 336.87 157.32 338.58 ;
   RECT 23.18 338.58 157.32 340.29 ;
   RECT 23.18 340.29 157.32 342.0 ;
   RECT 23.18 342.0 157.32 343.71 ;
   RECT 23.18 343.71 157.32 345.42 ;
   RECT 23.18 345.42 157.32 347.13 ;
   RECT 23.18 347.13 157.32 348.84 ;
   RECT 23.18 348.84 157.32 350.55 ;
   RECT 23.18 350.55 157.32 352.26 ;
   RECT 23.18 352.26 157.32 353.97 ;
   RECT 23.18 353.97 157.32 355.68 ;
   RECT 0.0 355.68 157.32 357.39 ;
   RECT 0.0 357.39 157.32 359.1 ;
   RECT 0.0 359.1 157.32 360.81 ;
   RECT 0.0 360.81 157.32 362.52 ;
   RECT 0.0 362.52 157.32 364.23 ;
   RECT 0.0 364.23 157.32 365.94 ;
   RECT 0.0 365.94 157.32 367.65 ;
   RECT 0.0 367.65 157.32 369.36 ;
   RECT 0.0 369.36 157.32 371.07 ;
   RECT 0.0 371.07 157.32 372.78 ;
   RECT 0.0 372.78 157.32 374.49 ;
   RECT 0.0 374.49 157.32 376.2 ;
   RECT 0.0 376.2 157.32 377.91 ;
   RECT 0.0 377.91 157.32 379.62 ;
   RECT 0.0 379.62 157.32 381.33 ;
   RECT 0.0 381.33 157.32 383.04 ;
   RECT 0.0 383.04 157.32 384.75 ;
   RECT 23.18 384.75 157.32 386.46 ;
   RECT 23.18 386.46 157.32 388.17 ;
   RECT 23.18 388.17 157.32 389.88 ;
   RECT 23.18 389.88 157.32 391.59 ;
   RECT 23.18 391.59 157.32 393.3 ;
   RECT 23.18 393.3 157.32 395.01 ;
   RECT 23.18 395.01 157.32 396.72 ;
   RECT 23.18 396.72 157.32 398.43 ;
   RECT 23.18 398.43 157.32 400.14 ;
   RECT 23.18 400.14 157.32 401.85 ;
   RECT 23.18 401.85 157.32 403.56 ;
   RECT 23.18 403.56 157.32 405.27 ;
   RECT 23.18 405.27 157.32 406.98 ;
   RECT 23.18 406.98 157.32 408.69 ;
   RECT 23.18 408.69 157.32 410.4 ;
   RECT 23.18 410.4 157.32 412.11 ;
   RECT 23.18 412.11 157.32 413.82 ;
   RECT 23.18 413.82 157.32 415.53 ;
   RECT 23.18 415.53 157.32 417.24 ;
   RECT 23.18 417.24 157.32 418.95 ;
   RECT 23.18 418.95 157.32 420.66 ;
   RECT 23.18 420.66 157.32 422.37 ;
   RECT 23.18 422.37 157.32 424.08 ;
   RECT 23.18 424.08 157.32 425.79 ;
   RECT 23.18 425.79 157.32 427.5 ;
   RECT 23.18 427.5 157.32 429.21 ;
   RECT 23.18 429.21 157.32 430.92 ;
   RECT 23.18 430.92 157.32 432.63 ;
   RECT 23.18 432.63 157.32 434.34 ;
   RECT 23.18 434.34 157.32 436.05 ;
   RECT 23.18 436.05 157.32 437.76 ;
   RECT 23.18 437.76 157.32 439.47 ;
   RECT 23.18 439.47 157.32 441.18 ;
   RECT 23.18 441.18 157.32 442.89 ;
   RECT 23.18 442.89 157.32 444.6 ;
   RECT 23.18 444.6 157.32 446.31 ;
   RECT 23.18 446.31 157.32 448.02 ;
   RECT 23.18 448.02 157.32 449.73 ;
   RECT 23.18 449.73 157.32 451.44 ;
   RECT 23.18 451.44 157.32 453.15 ;
   RECT 23.18 453.15 157.32 454.86 ;
   RECT 23.18 454.86 157.32 456.57 ;
   RECT 23.18 456.57 157.32 458.28 ;
   RECT 23.18 458.28 157.32 459.99 ;
   RECT 23.18 459.99 157.32 461.7 ;
   RECT 23.18 461.7 157.32 463.41 ;
   RECT 23.18 463.41 157.32 465.12 ;
   RECT 23.18 465.12 157.32 466.83 ;
   RECT 23.18 466.83 157.32 468.54 ;
   RECT 23.18 468.54 157.32 470.25 ;
   RECT 23.18 470.25 157.32 471.96 ;
   RECT 23.18 471.96 157.32 473.67 ;
   RECT 23.18 473.67 157.32 475.38 ;
   RECT 23.18 475.38 157.32 477.09 ;
   RECT 23.18 477.09 157.32 478.8 ;
   RECT 23.18 478.8 157.32 480.51 ;
   RECT 23.18 480.51 157.32 482.22 ;
   RECT 23.18 482.22 157.32 483.93 ;
   RECT 23.18 483.93 157.32 485.64 ;
   RECT 23.18 485.64 157.32 487.35 ;
   RECT 23.18 487.35 157.32 489.06 ;
   RECT 23.18 489.06 157.32 490.77 ;
   RECT 23.18 490.77 157.32 492.48 ;
   RECT 23.18 492.48 157.32 494.19 ;
   RECT 23.18 494.19 157.32 495.9 ;
   RECT 23.18 495.9 157.32 497.61 ;
   RECT 23.18 497.61 157.32 499.32 ;
   RECT 23.18 499.32 157.32 501.03 ;
   RECT 23.18 501.03 157.32 502.74 ;
   RECT 23.18 502.74 157.32 504.45 ;
   RECT 23.18 504.45 157.32 506.16 ;
   RECT 23.18 506.16 157.32 507.87 ;
   RECT 23.18 507.87 157.32 509.58 ;
   RECT 23.18 509.58 157.32 511.29 ;
   RECT 23.18 511.29 157.32 513.0 ;
   RECT 23.18 513.0 157.32 514.71 ;
   RECT 23.18 514.71 157.32 516.42 ;
   RECT 23.18 516.42 157.32 518.13 ;
   RECT 23.18 518.13 157.32 519.84 ;
   RECT 23.18 519.84 157.32 521.55 ;
   RECT 23.18 521.55 157.32 523.26 ;
   RECT 23.18 523.26 157.32 524.97 ;
   RECT 23.18 524.97 157.32 526.68 ;
   RECT 23.18 526.68 157.32 528.39 ;
   RECT 23.18 528.39 157.32 530.1 ;
   RECT 23.18 530.1 157.32 531.81 ;
   RECT 23.18 531.81 157.32 533.52 ;
   RECT 23.18 533.52 157.32 535.23 ;
   RECT 23.18 535.23 157.32 536.94 ;
   RECT 23.18 536.94 157.32 538.65 ;
   RECT 23.18 538.65 157.32 540.36 ;
   RECT 23.18 540.36 157.32 542.07 ;
   RECT 23.18 542.07 157.32 543.78 ;
   RECT 23.18 543.78 157.32 545.49 ;
   RECT 23.18 545.49 157.32 547.2 ;
   RECT 23.18 547.2 157.32 548.91 ;
   RECT 23.18 548.91 157.32 550.62 ;
   RECT 23.18 550.62 157.32 552.33 ;
   RECT 23.18 552.33 157.32 554.04 ;
   RECT 23.18 554.04 157.32 555.75 ;
   RECT 23.18 555.75 157.32 557.46 ;
   RECT 23.18 557.46 157.32 559.17 ;
   RECT 23.18 559.17 157.32 560.88 ;
   RECT 23.18 560.88 157.32 562.59 ;
   RECT 23.18 562.59 157.32 564.3 ;
   RECT 23.18 564.3 157.32 566.01 ;
   RECT 23.18 566.01 157.32 567.72 ;
   RECT 23.18 567.72 157.32 569.43 ;
   RECT 23.18 569.43 157.32 571.14 ;
   RECT 23.18 571.14 157.32 572.85 ;
   RECT 23.18 572.85 157.32 574.56 ;
   RECT 23.18 574.56 157.32 576.27 ;
   RECT 23.18 576.27 157.32 577.98 ;
   RECT 23.18 577.98 157.32 579.69 ;
   RECT 23.18 579.69 157.32 581.4 ;
   RECT 23.18 581.4 157.32 583.11 ;
   RECT 23.18 583.11 157.32 584.82 ;
   RECT 23.18 584.82 157.32 586.53 ;
   RECT 23.18 586.53 157.32 588.24 ;
   RECT 23.18 588.24 157.32 589.95 ;
   RECT 23.18 589.95 157.32 591.66 ;
   RECT 23.18 591.66 157.32 593.37 ;
   RECT 23.18 593.37 157.32 595.08 ;
   RECT 23.18 595.08 157.32 596.79 ;
   RECT 23.18 596.79 157.32 598.5 ;
   RECT 23.18 598.5 157.32 600.21 ;
   RECT 23.18 600.21 157.32 601.92 ;
   RECT 23.18 601.92 157.32 603.63 ;
   RECT 23.18 603.63 157.32 605.34 ;
   RECT 23.18 605.34 157.32 607.05 ;
   RECT 23.18 607.05 157.32 608.76 ;
   RECT 23.18 608.76 157.32 610.47 ;
   RECT 23.18 610.47 157.32 612.18 ;
   RECT 23.18 612.18 157.32 613.89 ;
   RECT 23.18 613.89 157.32 615.6 ;
   RECT 23.18 615.6 157.32 617.31 ;
   RECT 23.18 617.31 157.32 619.02 ;
   RECT 23.18 619.02 157.32 620.73 ;
   RECT 23.18 620.73 157.32 622.44 ;
   RECT 23.18 622.44 157.32 624.15 ;
   RECT 23.18 624.15 157.32 625.86 ;
   RECT 23.18 625.86 157.32 627.57 ;
   RECT 23.18 627.57 157.32 629.28 ;
   RECT 23.18 629.28 157.32 630.99 ;
   RECT 23.18 630.99 157.32 632.7 ;
   RECT 23.18 632.7 157.32 634.41 ;
   RECT 23.18 634.41 157.32 636.12 ;
   RECT 23.18 636.12 157.32 637.83 ;
   RECT 23.18 637.83 157.32 639.54 ;
   RECT 23.18 639.54 157.32 641.25 ;
   RECT 23.18 641.25 157.32 642.96 ;
   RECT 23.18 642.96 157.32 644.67 ;
   RECT 23.18 644.67 157.32 646.38 ;
   RECT 23.18 646.38 157.32 648.09 ;
   RECT 23.18 648.09 157.32 649.8 ;
   RECT 23.18 649.8 157.32 651.51 ;
   RECT 23.18 651.51 157.32 653.22 ;
   RECT 23.18 653.22 157.32 654.93 ;
   RECT 23.18 654.93 157.32 656.64 ;
   RECT 23.18 656.64 157.32 658.35 ;
   RECT 23.18 658.35 157.32 660.06 ;
   RECT 23.18 660.06 157.32 661.77 ;
   RECT 23.18 661.77 157.32 663.48 ;
   RECT 23.18 663.48 157.32 665.19 ;
   RECT 23.18 665.19 157.32 666.9 ;
   RECT 23.18 666.9 157.32 668.61 ;
   RECT 23.18 668.61 157.32 670.32 ;
   RECT 23.18 670.32 157.32 672.03 ;
   RECT 23.18 672.03 157.32 673.74 ;
   RECT 23.18 673.74 157.32 675.45 ;
   RECT 23.18 675.45 157.32 677.16 ;
   RECT 23.18 677.16 157.32 678.87 ;
   RECT 23.18 678.87 157.32 680.58 ;
   RECT 23.18 680.58 157.32 682.29 ;
   RECT 23.18 682.29 157.32 684.0 ;
   RECT 23.18 684.0 157.32 685.71 ;
   RECT 23.18 685.71 157.32 687.42 ;
   RECT 23.18 687.42 157.32 689.13 ;
   RECT 23.18 689.13 157.32 690.84 ;
   RECT 23.18 690.84 157.32 692.55 ;
   RECT 23.18 692.55 157.32 694.26 ;
   RECT 23.18 694.26 157.32 695.97 ;
   RECT 23.18 695.97 157.32 697.68 ;
   RECT 23.18 697.68 157.32 699.39 ;
   RECT 23.18 699.39 157.32 701.1 ;
   RECT 23.18 701.1 157.32 702.81 ;
   RECT 23.18 702.81 157.32 704.52 ;
   RECT 23.18 704.52 157.32 706.23 ;
   RECT 23.18 706.23 157.32 707.94 ;
   RECT 23.18 707.94 157.32 709.65 ;
   RECT 23.18 709.65 157.32 711.36 ;
   RECT 23.18 711.36 157.32 713.07 ;
   RECT 23.18 713.07 157.32 714.78 ;
   RECT 23.18 714.78 157.32 716.49 ;
   RECT 23.18 716.49 157.32 718.2 ;
   RECT 23.18 718.2 157.32 719.91 ;
   RECT 23.18 719.91 157.32 721.62 ;
   RECT 23.18 721.62 157.32 723.33 ;
   RECT 23.18 723.33 157.32 725.04 ;
   RECT 23.18 725.04 157.32 726.75 ;
   RECT 23.18 726.75 157.32 728.46 ;
   RECT 23.18 728.46 157.32 730.17 ;
   RECT 23.18 730.17 157.32 731.88 ;
   RECT 23.18 731.88 157.32 733.59 ;
   RECT 23.18 733.59 157.32 735.3 ;
   RECT 23.18 735.3 157.32 737.01 ;
   RECT 23.18 737.01 157.32 738.72 ;
   RECT 23.18 738.72 157.32 740.43 ;
   RECT 23.18 740.43 157.32 742.14 ;
   RECT 23.18 742.14 157.32 743.85 ;
   RECT 23.18 743.85 157.32 745.56 ;
   RECT 23.18 745.56 157.32 747.27 ;
   RECT 23.18 747.27 157.32 748.98 ;
   RECT 23.18 748.98 157.32 750.69 ;
   RECT 23.18 750.69 157.32 752.4 ;
   RECT 23.18 752.4 157.32 754.11 ;
  LAYER via1 ;
   RECT 23.18 0.0 157.32 1.71 ;
   RECT 23.18 1.71 157.32 3.42 ;
   RECT 23.18 3.42 157.32 5.13 ;
   RECT 23.18 5.13 157.32 6.84 ;
   RECT 23.18 6.84 157.32 8.55 ;
   RECT 23.18 8.55 157.32 10.26 ;
   RECT 23.18 10.26 157.32 11.97 ;
   RECT 23.18 11.97 157.32 13.68 ;
   RECT 23.18 13.68 157.32 15.39 ;
   RECT 23.18 15.39 157.32 17.1 ;
   RECT 23.18 17.1 157.32 18.81 ;
   RECT 23.18 18.81 157.32 20.52 ;
   RECT 23.18 20.52 157.32 22.23 ;
   RECT 23.18 22.23 157.32 23.94 ;
   RECT 23.18 23.94 157.32 25.65 ;
   RECT 23.18 25.65 157.32 27.36 ;
   RECT 23.18 27.36 157.32 29.07 ;
   RECT 23.18 29.07 157.32 30.78 ;
   RECT 23.18 30.78 157.32 32.49 ;
   RECT 23.18 32.49 157.32 34.2 ;
   RECT 23.18 34.2 157.32 35.91 ;
   RECT 23.18 35.91 157.32 37.62 ;
   RECT 23.18 37.62 157.32 39.33 ;
   RECT 23.18 39.33 157.32 41.04 ;
   RECT 23.18 41.04 157.32 42.75 ;
   RECT 23.18 42.75 157.32 44.46 ;
   RECT 23.18 44.46 157.32 46.17 ;
   RECT 23.18 46.17 157.32 47.88 ;
   RECT 23.18 47.88 157.32 49.59 ;
   RECT 23.18 49.59 157.32 51.3 ;
   RECT 23.18 51.3 157.32 53.01 ;
   RECT 23.18 53.01 157.32 54.72 ;
   RECT 23.18 54.72 157.32 56.43 ;
   RECT 23.18 56.43 157.32 58.14 ;
   RECT 23.18 58.14 157.32 59.85 ;
   RECT 23.18 59.85 157.32 61.56 ;
   RECT 23.18 61.56 157.32 63.27 ;
   RECT 23.18 63.27 157.32 64.98 ;
   RECT 23.18 64.98 157.32 66.69 ;
   RECT 23.18 66.69 157.32 68.4 ;
   RECT 23.18 68.4 157.32 70.11 ;
   RECT 23.18 70.11 157.32 71.82 ;
   RECT 23.18 71.82 157.32 73.53 ;
   RECT 23.18 73.53 157.32 75.24 ;
   RECT 23.18 75.24 157.32 76.95 ;
   RECT 23.18 76.95 157.32 78.66 ;
   RECT 23.18 78.66 157.32 80.37 ;
   RECT 23.18 80.37 157.32 82.08 ;
   RECT 23.18 82.08 157.32 83.79 ;
   RECT 23.18 83.79 157.32 85.5 ;
   RECT 23.18 85.5 157.32 87.21 ;
   RECT 23.18 87.21 157.32 88.92 ;
   RECT 23.18 88.92 157.32 90.63 ;
   RECT 23.18 90.63 157.32 92.34 ;
   RECT 23.18 92.34 157.32 94.05 ;
   RECT 23.18 94.05 157.32 95.76 ;
   RECT 23.18 95.76 157.32 97.47 ;
   RECT 23.18 97.47 157.32 99.18 ;
   RECT 23.18 99.18 157.32 100.89 ;
   RECT 23.18 100.89 157.32 102.6 ;
   RECT 23.18 102.6 157.32 104.31 ;
   RECT 23.18 104.31 157.32 106.02 ;
   RECT 23.18 106.02 157.32 107.73 ;
   RECT 23.18 107.73 157.32 109.44 ;
   RECT 23.18 109.44 157.32 111.15 ;
   RECT 23.18 111.15 157.32 112.86 ;
   RECT 23.18 112.86 157.32 114.57 ;
   RECT 23.18 114.57 157.32 116.28 ;
   RECT 23.18 116.28 157.32 117.99 ;
   RECT 23.18 117.99 157.32 119.7 ;
   RECT 23.18 119.7 157.32 121.41 ;
   RECT 23.18 121.41 157.32 123.12 ;
   RECT 23.18 123.12 157.32 124.83 ;
   RECT 23.18 124.83 157.32 126.54 ;
   RECT 23.18 126.54 157.32 128.25 ;
   RECT 23.18 128.25 157.32 129.96 ;
   RECT 23.18 129.96 157.32 131.67 ;
   RECT 23.18 131.67 157.32 133.38 ;
   RECT 23.18 133.38 157.32 135.09 ;
   RECT 23.18 135.09 157.32 136.8 ;
   RECT 23.18 136.8 157.32 138.51 ;
   RECT 23.18 138.51 157.32 140.22 ;
   RECT 23.18 140.22 157.32 141.93 ;
   RECT 23.18 141.93 157.32 143.64 ;
   RECT 23.18 143.64 157.32 145.35 ;
   RECT 23.18 145.35 157.32 147.06 ;
   RECT 23.18 147.06 157.32 148.77 ;
   RECT 23.18 148.77 157.32 150.48 ;
   RECT 23.18 150.48 157.32 152.19 ;
   RECT 23.18 152.19 157.32 153.9 ;
   RECT 23.18 153.9 157.32 155.61 ;
   RECT 23.18 155.61 157.32 157.32 ;
   RECT 23.18 157.32 157.32 159.03 ;
   RECT 23.18 159.03 157.32 160.74 ;
   RECT 23.18 160.74 157.32 162.45 ;
   RECT 23.18 162.45 157.32 164.16 ;
   RECT 23.18 164.16 157.32 165.87 ;
   RECT 23.18 165.87 157.32 167.58 ;
   RECT 23.18 167.58 157.32 169.29 ;
   RECT 23.18 169.29 157.32 171.0 ;
   RECT 23.18 171.0 157.32 172.71 ;
   RECT 23.18 172.71 157.32 174.42 ;
   RECT 23.18 174.42 157.32 176.13 ;
   RECT 23.18 176.13 157.32 177.84 ;
   RECT 23.18 177.84 157.32 179.55 ;
   RECT 23.18 179.55 157.32 181.26 ;
   RECT 23.18 181.26 157.32 182.97 ;
   RECT 23.18 182.97 157.32 184.68 ;
   RECT 23.18 184.68 157.32 186.39 ;
   RECT 23.18 186.39 157.32 188.1 ;
   RECT 23.18 188.1 157.32 189.81 ;
   RECT 23.18 189.81 157.32 191.52 ;
   RECT 23.18 191.52 157.32 193.23 ;
   RECT 23.18 193.23 157.32 194.94 ;
   RECT 23.18 194.94 157.32 196.65 ;
   RECT 23.18 196.65 157.32 198.36 ;
   RECT 23.18 198.36 157.32 200.07 ;
   RECT 23.18 200.07 157.32 201.78 ;
   RECT 23.18 201.78 157.32 203.49 ;
   RECT 23.18 203.49 157.32 205.2 ;
   RECT 23.18 205.2 157.32 206.91 ;
   RECT 23.18 206.91 157.32 208.62 ;
   RECT 23.18 208.62 157.32 210.33 ;
   RECT 23.18 210.33 157.32 212.04 ;
   RECT 23.18 212.04 157.32 213.75 ;
   RECT 23.18 213.75 157.32 215.46 ;
   RECT 23.18 215.46 157.32 217.17 ;
   RECT 23.18 217.17 157.32 218.88 ;
   RECT 23.18 218.88 157.32 220.59 ;
   RECT 23.18 220.59 157.32 222.3 ;
   RECT 23.18 222.3 157.32 224.01 ;
   RECT 23.18 224.01 157.32 225.72 ;
   RECT 23.18 225.72 157.32 227.43 ;
   RECT 23.18 227.43 157.32 229.14 ;
   RECT 23.18 229.14 157.32 230.85 ;
   RECT 23.18 230.85 157.32 232.56 ;
   RECT 23.18 232.56 157.32 234.27 ;
   RECT 23.18 234.27 157.32 235.98 ;
   RECT 23.18 235.98 157.32 237.69 ;
   RECT 23.18 237.69 157.32 239.4 ;
   RECT 23.18 239.4 157.32 241.11 ;
   RECT 23.18 241.11 157.32 242.82 ;
   RECT 23.18 242.82 157.32 244.53 ;
   RECT 23.18 244.53 157.32 246.24 ;
   RECT 23.18 246.24 157.32 247.95 ;
   RECT 23.18 247.95 157.32 249.66 ;
   RECT 23.18 249.66 157.32 251.37 ;
   RECT 23.18 251.37 157.32 253.08 ;
   RECT 23.18 253.08 157.32 254.79 ;
   RECT 23.18 254.79 157.32 256.5 ;
   RECT 23.18 256.5 157.32 258.21 ;
   RECT 23.18 258.21 157.32 259.92 ;
   RECT 23.18 259.92 157.32 261.63 ;
   RECT 23.18 261.63 157.32 263.34 ;
   RECT 23.18 263.34 157.32 265.05 ;
   RECT 23.18 265.05 157.32 266.76 ;
   RECT 23.18 266.76 157.32 268.47 ;
   RECT 23.18 268.47 157.32 270.18 ;
   RECT 23.18 270.18 157.32 271.89 ;
   RECT 23.18 271.89 157.32 273.6 ;
   RECT 23.18 273.6 157.32 275.31 ;
   RECT 23.18 275.31 157.32 277.02 ;
   RECT 23.18 277.02 157.32 278.73 ;
   RECT 23.18 278.73 157.32 280.44 ;
   RECT 23.18 280.44 157.32 282.15 ;
   RECT 23.18 282.15 157.32 283.86 ;
   RECT 23.18 283.86 157.32 285.57 ;
   RECT 23.18 285.57 157.32 287.28 ;
   RECT 23.18 287.28 157.32 288.99 ;
   RECT 23.18 288.99 157.32 290.7 ;
   RECT 23.18 290.7 157.32 292.41 ;
   RECT 23.18 292.41 157.32 294.12 ;
   RECT 23.18 294.12 157.32 295.83 ;
   RECT 23.18 295.83 157.32 297.54 ;
   RECT 23.18 297.54 157.32 299.25 ;
   RECT 23.18 299.25 157.32 300.96 ;
   RECT 23.18 300.96 157.32 302.67 ;
   RECT 23.18 302.67 157.32 304.38 ;
   RECT 23.18 304.38 157.32 306.09 ;
   RECT 23.18 306.09 157.32 307.8 ;
   RECT 23.18 307.8 157.32 309.51 ;
   RECT 23.18 309.51 157.32 311.22 ;
   RECT 23.18 311.22 157.32 312.93 ;
   RECT 23.18 312.93 157.32 314.64 ;
   RECT 23.18 314.64 157.32 316.35 ;
   RECT 23.18 316.35 157.32 318.06 ;
   RECT 23.18 318.06 157.32 319.77 ;
   RECT 23.18 319.77 157.32 321.48 ;
   RECT 23.18 321.48 157.32 323.19 ;
   RECT 23.18 323.19 157.32 324.9 ;
   RECT 23.18 324.9 157.32 326.61 ;
   RECT 23.18 326.61 157.32 328.32 ;
   RECT 23.18 328.32 157.32 330.03 ;
   RECT 23.18 330.03 157.32 331.74 ;
   RECT 23.18 331.74 157.32 333.45 ;
   RECT 23.18 333.45 157.32 335.16 ;
   RECT 23.18 335.16 157.32 336.87 ;
   RECT 23.18 336.87 157.32 338.58 ;
   RECT 23.18 338.58 157.32 340.29 ;
   RECT 23.18 340.29 157.32 342.0 ;
   RECT 23.18 342.0 157.32 343.71 ;
   RECT 23.18 343.71 157.32 345.42 ;
   RECT 23.18 345.42 157.32 347.13 ;
   RECT 23.18 347.13 157.32 348.84 ;
   RECT 23.18 348.84 157.32 350.55 ;
   RECT 23.18 350.55 157.32 352.26 ;
   RECT 23.18 352.26 157.32 353.97 ;
   RECT 23.18 353.97 157.32 355.68 ;
   RECT 0.0 355.68 157.32 357.39 ;
   RECT 0.0 357.39 157.32 359.1 ;
   RECT 0.0 359.1 157.32 360.81 ;
   RECT 0.0 360.81 157.32 362.52 ;
   RECT 0.0 362.52 157.32 364.23 ;
   RECT 0.0 364.23 157.32 365.94 ;
   RECT 0.0 365.94 157.32 367.65 ;
   RECT 0.0 367.65 157.32 369.36 ;
   RECT 0.0 369.36 157.32 371.07 ;
   RECT 0.0 371.07 157.32 372.78 ;
   RECT 0.0 372.78 157.32 374.49 ;
   RECT 0.0 374.49 157.32 376.2 ;
   RECT 0.0 376.2 157.32 377.91 ;
   RECT 0.0 377.91 157.32 379.62 ;
   RECT 0.0 379.62 157.32 381.33 ;
   RECT 0.0 381.33 157.32 383.04 ;
   RECT 0.0 383.04 157.32 384.75 ;
   RECT 23.18 384.75 157.32 386.46 ;
   RECT 23.18 386.46 157.32 388.17 ;
   RECT 23.18 388.17 157.32 389.88 ;
   RECT 23.18 389.88 157.32 391.59 ;
   RECT 23.18 391.59 157.32 393.3 ;
   RECT 23.18 393.3 157.32 395.01 ;
   RECT 23.18 395.01 157.32 396.72 ;
   RECT 23.18 396.72 157.32 398.43 ;
   RECT 23.18 398.43 157.32 400.14 ;
   RECT 23.18 400.14 157.32 401.85 ;
   RECT 23.18 401.85 157.32 403.56 ;
   RECT 23.18 403.56 157.32 405.27 ;
   RECT 23.18 405.27 157.32 406.98 ;
   RECT 23.18 406.98 157.32 408.69 ;
   RECT 23.18 408.69 157.32 410.4 ;
   RECT 23.18 410.4 157.32 412.11 ;
   RECT 23.18 412.11 157.32 413.82 ;
   RECT 23.18 413.82 157.32 415.53 ;
   RECT 23.18 415.53 157.32 417.24 ;
   RECT 23.18 417.24 157.32 418.95 ;
   RECT 23.18 418.95 157.32 420.66 ;
   RECT 23.18 420.66 157.32 422.37 ;
   RECT 23.18 422.37 157.32 424.08 ;
   RECT 23.18 424.08 157.32 425.79 ;
   RECT 23.18 425.79 157.32 427.5 ;
   RECT 23.18 427.5 157.32 429.21 ;
   RECT 23.18 429.21 157.32 430.92 ;
   RECT 23.18 430.92 157.32 432.63 ;
   RECT 23.18 432.63 157.32 434.34 ;
   RECT 23.18 434.34 157.32 436.05 ;
   RECT 23.18 436.05 157.32 437.76 ;
   RECT 23.18 437.76 157.32 439.47 ;
   RECT 23.18 439.47 157.32 441.18 ;
   RECT 23.18 441.18 157.32 442.89 ;
   RECT 23.18 442.89 157.32 444.6 ;
   RECT 23.18 444.6 157.32 446.31 ;
   RECT 23.18 446.31 157.32 448.02 ;
   RECT 23.18 448.02 157.32 449.73 ;
   RECT 23.18 449.73 157.32 451.44 ;
   RECT 23.18 451.44 157.32 453.15 ;
   RECT 23.18 453.15 157.32 454.86 ;
   RECT 23.18 454.86 157.32 456.57 ;
   RECT 23.18 456.57 157.32 458.28 ;
   RECT 23.18 458.28 157.32 459.99 ;
   RECT 23.18 459.99 157.32 461.7 ;
   RECT 23.18 461.7 157.32 463.41 ;
   RECT 23.18 463.41 157.32 465.12 ;
   RECT 23.18 465.12 157.32 466.83 ;
   RECT 23.18 466.83 157.32 468.54 ;
   RECT 23.18 468.54 157.32 470.25 ;
   RECT 23.18 470.25 157.32 471.96 ;
   RECT 23.18 471.96 157.32 473.67 ;
   RECT 23.18 473.67 157.32 475.38 ;
   RECT 23.18 475.38 157.32 477.09 ;
   RECT 23.18 477.09 157.32 478.8 ;
   RECT 23.18 478.8 157.32 480.51 ;
   RECT 23.18 480.51 157.32 482.22 ;
   RECT 23.18 482.22 157.32 483.93 ;
   RECT 23.18 483.93 157.32 485.64 ;
   RECT 23.18 485.64 157.32 487.35 ;
   RECT 23.18 487.35 157.32 489.06 ;
   RECT 23.18 489.06 157.32 490.77 ;
   RECT 23.18 490.77 157.32 492.48 ;
   RECT 23.18 492.48 157.32 494.19 ;
   RECT 23.18 494.19 157.32 495.9 ;
   RECT 23.18 495.9 157.32 497.61 ;
   RECT 23.18 497.61 157.32 499.32 ;
   RECT 23.18 499.32 157.32 501.03 ;
   RECT 23.18 501.03 157.32 502.74 ;
   RECT 23.18 502.74 157.32 504.45 ;
   RECT 23.18 504.45 157.32 506.16 ;
   RECT 23.18 506.16 157.32 507.87 ;
   RECT 23.18 507.87 157.32 509.58 ;
   RECT 23.18 509.58 157.32 511.29 ;
   RECT 23.18 511.29 157.32 513.0 ;
   RECT 23.18 513.0 157.32 514.71 ;
   RECT 23.18 514.71 157.32 516.42 ;
   RECT 23.18 516.42 157.32 518.13 ;
   RECT 23.18 518.13 157.32 519.84 ;
   RECT 23.18 519.84 157.32 521.55 ;
   RECT 23.18 521.55 157.32 523.26 ;
   RECT 23.18 523.26 157.32 524.97 ;
   RECT 23.18 524.97 157.32 526.68 ;
   RECT 23.18 526.68 157.32 528.39 ;
   RECT 23.18 528.39 157.32 530.1 ;
   RECT 23.18 530.1 157.32 531.81 ;
   RECT 23.18 531.81 157.32 533.52 ;
   RECT 23.18 533.52 157.32 535.23 ;
   RECT 23.18 535.23 157.32 536.94 ;
   RECT 23.18 536.94 157.32 538.65 ;
   RECT 23.18 538.65 157.32 540.36 ;
   RECT 23.18 540.36 157.32 542.07 ;
   RECT 23.18 542.07 157.32 543.78 ;
   RECT 23.18 543.78 157.32 545.49 ;
   RECT 23.18 545.49 157.32 547.2 ;
   RECT 23.18 547.2 157.32 548.91 ;
   RECT 23.18 548.91 157.32 550.62 ;
   RECT 23.18 550.62 157.32 552.33 ;
   RECT 23.18 552.33 157.32 554.04 ;
   RECT 23.18 554.04 157.32 555.75 ;
   RECT 23.18 555.75 157.32 557.46 ;
   RECT 23.18 557.46 157.32 559.17 ;
   RECT 23.18 559.17 157.32 560.88 ;
   RECT 23.18 560.88 157.32 562.59 ;
   RECT 23.18 562.59 157.32 564.3 ;
   RECT 23.18 564.3 157.32 566.01 ;
   RECT 23.18 566.01 157.32 567.72 ;
   RECT 23.18 567.72 157.32 569.43 ;
   RECT 23.18 569.43 157.32 571.14 ;
   RECT 23.18 571.14 157.32 572.85 ;
   RECT 23.18 572.85 157.32 574.56 ;
   RECT 23.18 574.56 157.32 576.27 ;
   RECT 23.18 576.27 157.32 577.98 ;
   RECT 23.18 577.98 157.32 579.69 ;
   RECT 23.18 579.69 157.32 581.4 ;
   RECT 23.18 581.4 157.32 583.11 ;
   RECT 23.18 583.11 157.32 584.82 ;
   RECT 23.18 584.82 157.32 586.53 ;
   RECT 23.18 586.53 157.32 588.24 ;
   RECT 23.18 588.24 157.32 589.95 ;
   RECT 23.18 589.95 157.32 591.66 ;
   RECT 23.18 591.66 157.32 593.37 ;
   RECT 23.18 593.37 157.32 595.08 ;
   RECT 23.18 595.08 157.32 596.79 ;
   RECT 23.18 596.79 157.32 598.5 ;
   RECT 23.18 598.5 157.32 600.21 ;
   RECT 23.18 600.21 157.32 601.92 ;
   RECT 23.18 601.92 157.32 603.63 ;
   RECT 23.18 603.63 157.32 605.34 ;
   RECT 23.18 605.34 157.32 607.05 ;
   RECT 23.18 607.05 157.32 608.76 ;
   RECT 23.18 608.76 157.32 610.47 ;
   RECT 23.18 610.47 157.32 612.18 ;
   RECT 23.18 612.18 157.32 613.89 ;
   RECT 23.18 613.89 157.32 615.6 ;
   RECT 23.18 615.6 157.32 617.31 ;
   RECT 23.18 617.31 157.32 619.02 ;
   RECT 23.18 619.02 157.32 620.73 ;
   RECT 23.18 620.73 157.32 622.44 ;
   RECT 23.18 622.44 157.32 624.15 ;
   RECT 23.18 624.15 157.32 625.86 ;
   RECT 23.18 625.86 157.32 627.57 ;
   RECT 23.18 627.57 157.32 629.28 ;
   RECT 23.18 629.28 157.32 630.99 ;
   RECT 23.18 630.99 157.32 632.7 ;
   RECT 23.18 632.7 157.32 634.41 ;
   RECT 23.18 634.41 157.32 636.12 ;
   RECT 23.18 636.12 157.32 637.83 ;
   RECT 23.18 637.83 157.32 639.54 ;
   RECT 23.18 639.54 157.32 641.25 ;
   RECT 23.18 641.25 157.32 642.96 ;
   RECT 23.18 642.96 157.32 644.67 ;
   RECT 23.18 644.67 157.32 646.38 ;
   RECT 23.18 646.38 157.32 648.09 ;
   RECT 23.18 648.09 157.32 649.8 ;
   RECT 23.18 649.8 157.32 651.51 ;
   RECT 23.18 651.51 157.32 653.22 ;
   RECT 23.18 653.22 157.32 654.93 ;
   RECT 23.18 654.93 157.32 656.64 ;
   RECT 23.18 656.64 157.32 658.35 ;
   RECT 23.18 658.35 157.32 660.06 ;
   RECT 23.18 660.06 157.32 661.77 ;
   RECT 23.18 661.77 157.32 663.48 ;
   RECT 23.18 663.48 157.32 665.19 ;
   RECT 23.18 665.19 157.32 666.9 ;
   RECT 23.18 666.9 157.32 668.61 ;
   RECT 23.18 668.61 157.32 670.32 ;
   RECT 23.18 670.32 157.32 672.03 ;
   RECT 23.18 672.03 157.32 673.74 ;
   RECT 23.18 673.74 157.32 675.45 ;
   RECT 23.18 675.45 157.32 677.16 ;
   RECT 23.18 677.16 157.32 678.87 ;
   RECT 23.18 678.87 157.32 680.58 ;
   RECT 23.18 680.58 157.32 682.29 ;
   RECT 23.18 682.29 157.32 684.0 ;
   RECT 23.18 684.0 157.32 685.71 ;
   RECT 23.18 685.71 157.32 687.42 ;
   RECT 23.18 687.42 157.32 689.13 ;
   RECT 23.18 689.13 157.32 690.84 ;
   RECT 23.18 690.84 157.32 692.55 ;
   RECT 23.18 692.55 157.32 694.26 ;
   RECT 23.18 694.26 157.32 695.97 ;
   RECT 23.18 695.97 157.32 697.68 ;
   RECT 23.18 697.68 157.32 699.39 ;
   RECT 23.18 699.39 157.32 701.1 ;
   RECT 23.18 701.1 157.32 702.81 ;
   RECT 23.18 702.81 157.32 704.52 ;
   RECT 23.18 704.52 157.32 706.23 ;
   RECT 23.18 706.23 157.32 707.94 ;
   RECT 23.18 707.94 157.32 709.65 ;
   RECT 23.18 709.65 157.32 711.36 ;
   RECT 23.18 711.36 157.32 713.07 ;
   RECT 23.18 713.07 157.32 714.78 ;
   RECT 23.18 714.78 157.32 716.49 ;
   RECT 23.18 716.49 157.32 718.2 ;
   RECT 23.18 718.2 157.32 719.91 ;
   RECT 23.18 719.91 157.32 721.62 ;
   RECT 23.18 721.62 157.32 723.33 ;
   RECT 23.18 723.33 157.32 725.04 ;
   RECT 23.18 725.04 157.32 726.75 ;
   RECT 23.18 726.75 157.32 728.46 ;
   RECT 23.18 728.46 157.32 730.17 ;
   RECT 23.18 730.17 157.32 731.88 ;
   RECT 23.18 731.88 157.32 733.59 ;
   RECT 23.18 733.59 157.32 735.3 ;
   RECT 23.18 735.3 157.32 737.01 ;
   RECT 23.18 737.01 157.32 738.72 ;
   RECT 23.18 738.72 157.32 740.43 ;
   RECT 23.18 740.43 157.32 742.14 ;
   RECT 23.18 742.14 157.32 743.85 ;
   RECT 23.18 743.85 157.32 745.56 ;
   RECT 23.18 745.56 157.32 747.27 ;
   RECT 23.18 747.27 157.32 748.98 ;
   RECT 23.18 748.98 157.32 750.69 ;
   RECT 23.18 750.69 157.32 752.4 ;
   RECT 23.18 752.4 157.32 754.11 ;
  LAYER metal2 ;
   RECT 23.18 0.0 157.32 1.71 ;
   RECT 23.18 1.71 157.32 3.42 ;
   RECT 23.18 3.42 157.32 5.13 ;
   RECT 23.18 5.13 157.32 6.84 ;
   RECT 23.18 6.84 157.32 8.55 ;
   RECT 23.18 8.55 157.32 10.26 ;
   RECT 23.18 10.26 157.32 11.97 ;
   RECT 23.18 11.97 157.32 13.68 ;
   RECT 23.18 13.68 157.32 15.39 ;
   RECT 23.18 15.39 157.32 17.1 ;
   RECT 23.18 17.1 157.32 18.81 ;
   RECT 23.18 18.81 157.32 20.52 ;
   RECT 23.18 20.52 157.32 22.23 ;
   RECT 23.18 22.23 157.32 23.94 ;
   RECT 23.18 23.94 157.32 25.65 ;
   RECT 23.18 25.65 157.32 27.36 ;
   RECT 23.18 27.36 157.32 29.07 ;
   RECT 23.18 29.07 157.32 30.78 ;
   RECT 23.18 30.78 157.32 32.49 ;
   RECT 23.18 32.49 157.32 34.2 ;
   RECT 23.18 34.2 157.32 35.91 ;
   RECT 23.18 35.91 157.32 37.62 ;
   RECT 23.18 37.62 157.32 39.33 ;
   RECT 23.18 39.33 157.32 41.04 ;
   RECT 23.18 41.04 157.32 42.75 ;
   RECT 23.18 42.75 157.32 44.46 ;
   RECT 23.18 44.46 157.32 46.17 ;
   RECT 23.18 46.17 157.32 47.88 ;
   RECT 23.18 47.88 157.32 49.59 ;
   RECT 23.18 49.59 157.32 51.3 ;
   RECT 23.18 51.3 157.32 53.01 ;
   RECT 23.18 53.01 157.32 54.72 ;
   RECT 23.18 54.72 157.32 56.43 ;
   RECT 23.18 56.43 157.32 58.14 ;
   RECT 23.18 58.14 157.32 59.85 ;
   RECT 23.18 59.85 157.32 61.56 ;
   RECT 23.18 61.56 157.32 63.27 ;
   RECT 23.18 63.27 157.32 64.98 ;
   RECT 23.18 64.98 157.32 66.69 ;
   RECT 23.18 66.69 157.32 68.4 ;
   RECT 23.18 68.4 157.32 70.11 ;
   RECT 23.18 70.11 157.32 71.82 ;
   RECT 23.18 71.82 157.32 73.53 ;
   RECT 23.18 73.53 157.32 75.24 ;
   RECT 23.18 75.24 157.32 76.95 ;
   RECT 23.18 76.95 157.32 78.66 ;
   RECT 23.18 78.66 157.32 80.37 ;
   RECT 23.18 80.37 157.32 82.08 ;
   RECT 23.18 82.08 157.32 83.79 ;
   RECT 23.18 83.79 157.32 85.5 ;
   RECT 23.18 85.5 157.32 87.21 ;
   RECT 23.18 87.21 157.32 88.92 ;
   RECT 23.18 88.92 157.32 90.63 ;
   RECT 23.18 90.63 157.32 92.34 ;
   RECT 23.18 92.34 157.32 94.05 ;
   RECT 23.18 94.05 157.32 95.76 ;
   RECT 23.18 95.76 157.32 97.47 ;
   RECT 23.18 97.47 157.32 99.18 ;
   RECT 23.18 99.18 157.32 100.89 ;
   RECT 23.18 100.89 157.32 102.6 ;
   RECT 23.18 102.6 157.32 104.31 ;
   RECT 23.18 104.31 157.32 106.02 ;
   RECT 23.18 106.02 157.32 107.73 ;
   RECT 23.18 107.73 157.32 109.44 ;
   RECT 23.18 109.44 157.32 111.15 ;
   RECT 23.18 111.15 157.32 112.86 ;
   RECT 23.18 112.86 157.32 114.57 ;
   RECT 23.18 114.57 157.32 116.28 ;
   RECT 23.18 116.28 157.32 117.99 ;
   RECT 23.18 117.99 157.32 119.7 ;
   RECT 23.18 119.7 157.32 121.41 ;
   RECT 23.18 121.41 157.32 123.12 ;
   RECT 23.18 123.12 157.32 124.83 ;
   RECT 23.18 124.83 157.32 126.54 ;
   RECT 23.18 126.54 157.32 128.25 ;
   RECT 23.18 128.25 157.32 129.96 ;
   RECT 23.18 129.96 157.32 131.67 ;
   RECT 23.18 131.67 157.32 133.38 ;
   RECT 23.18 133.38 157.32 135.09 ;
   RECT 23.18 135.09 157.32 136.8 ;
   RECT 23.18 136.8 157.32 138.51 ;
   RECT 23.18 138.51 157.32 140.22 ;
   RECT 23.18 140.22 157.32 141.93 ;
   RECT 23.18 141.93 157.32 143.64 ;
   RECT 23.18 143.64 157.32 145.35 ;
   RECT 23.18 145.35 157.32 147.06 ;
   RECT 23.18 147.06 157.32 148.77 ;
   RECT 23.18 148.77 157.32 150.48 ;
   RECT 23.18 150.48 157.32 152.19 ;
   RECT 23.18 152.19 157.32 153.9 ;
   RECT 23.18 153.9 157.32 155.61 ;
   RECT 23.18 155.61 157.32 157.32 ;
   RECT 23.18 157.32 157.32 159.03 ;
   RECT 23.18 159.03 157.32 160.74 ;
   RECT 23.18 160.74 157.32 162.45 ;
   RECT 23.18 162.45 157.32 164.16 ;
   RECT 23.18 164.16 157.32 165.87 ;
   RECT 23.18 165.87 157.32 167.58 ;
   RECT 23.18 167.58 157.32 169.29 ;
   RECT 23.18 169.29 157.32 171.0 ;
   RECT 23.18 171.0 157.32 172.71 ;
   RECT 23.18 172.71 157.32 174.42 ;
   RECT 23.18 174.42 157.32 176.13 ;
   RECT 23.18 176.13 157.32 177.84 ;
   RECT 23.18 177.84 157.32 179.55 ;
   RECT 23.18 179.55 157.32 181.26 ;
   RECT 23.18 181.26 157.32 182.97 ;
   RECT 23.18 182.97 157.32 184.68 ;
   RECT 23.18 184.68 157.32 186.39 ;
   RECT 23.18 186.39 157.32 188.1 ;
   RECT 23.18 188.1 157.32 189.81 ;
   RECT 23.18 189.81 157.32 191.52 ;
   RECT 23.18 191.52 157.32 193.23 ;
   RECT 23.18 193.23 157.32 194.94 ;
   RECT 23.18 194.94 157.32 196.65 ;
   RECT 23.18 196.65 157.32 198.36 ;
   RECT 23.18 198.36 157.32 200.07 ;
   RECT 23.18 200.07 157.32 201.78 ;
   RECT 23.18 201.78 157.32 203.49 ;
   RECT 23.18 203.49 157.32 205.2 ;
   RECT 23.18 205.2 157.32 206.91 ;
   RECT 23.18 206.91 157.32 208.62 ;
   RECT 23.18 208.62 157.32 210.33 ;
   RECT 23.18 210.33 157.32 212.04 ;
   RECT 23.18 212.04 157.32 213.75 ;
   RECT 23.18 213.75 157.32 215.46 ;
   RECT 23.18 215.46 157.32 217.17 ;
   RECT 23.18 217.17 157.32 218.88 ;
   RECT 23.18 218.88 157.32 220.59 ;
   RECT 23.18 220.59 157.32 222.3 ;
   RECT 23.18 222.3 157.32 224.01 ;
   RECT 23.18 224.01 157.32 225.72 ;
   RECT 23.18 225.72 157.32 227.43 ;
   RECT 23.18 227.43 157.32 229.14 ;
   RECT 23.18 229.14 157.32 230.85 ;
   RECT 23.18 230.85 157.32 232.56 ;
   RECT 23.18 232.56 157.32 234.27 ;
   RECT 23.18 234.27 157.32 235.98 ;
   RECT 23.18 235.98 157.32 237.69 ;
   RECT 23.18 237.69 157.32 239.4 ;
   RECT 23.18 239.4 157.32 241.11 ;
   RECT 23.18 241.11 157.32 242.82 ;
   RECT 23.18 242.82 157.32 244.53 ;
   RECT 23.18 244.53 157.32 246.24 ;
   RECT 23.18 246.24 157.32 247.95 ;
   RECT 23.18 247.95 157.32 249.66 ;
   RECT 23.18 249.66 157.32 251.37 ;
   RECT 23.18 251.37 157.32 253.08 ;
   RECT 23.18 253.08 157.32 254.79 ;
   RECT 23.18 254.79 157.32 256.5 ;
   RECT 23.18 256.5 157.32 258.21 ;
   RECT 23.18 258.21 157.32 259.92 ;
   RECT 23.18 259.92 157.32 261.63 ;
   RECT 23.18 261.63 157.32 263.34 ;
   RECT 23.18 263.34 157.32 265.05 ;
   RECT 23.18 265.05 157.32 266.76 ;
   RECT 23.18 266.76 157.32 268.47 ;
   RECT 23.18 268.47 157.32 270.18 ;
   RECT 23.18 270.18 157.32 271.89 ;
   RECT 23.18 271.89 157.32 273.6 ;
   RECT 23.18 273.6 157.32 275.31 ;
   RECT 23.18 275.31 157.32 277.02 ;
   RECT 23.18 277.02 157.32 278.73 ;
   RECT 23.18 278.73 157.32 280.44 ;
   RECT 23.18 280.44 157.32 282.15 ;
   RECT 23.18 282.15 157.32 283.86 ;
   RECT 23.18 283.86 157.32 285.57 ;
   RECT 23.18 285.57 157.32 287.28 ;
   RECT 23.18 287.28 157.32 288.99 ;
   RECT 23.18 288.99 157.32 290.7 ;
   RECT 23.18 290.7 157.32 292.41 ;
   RECT 23.18 292.41 157.32 294.12 ;
   RECT 23.18 294.12 157.32 295.83 ;
   RECT 23.18 295.83 157.32 297.54 ;
   RECT 23.18 297.54 157.32 299.25 ;
   RECT 23.18 299.25 157.32 300.96 ;
   RECT 23.18 300.96 157.32 302.67 ;
   RECT 23.18 302.67 157.32 304.38 ;
   RECT 23.18 304.38 157.32 306.09 ;
   RECT 23.18 306.09 157.32 307.8 ;
   RECT 23.18 307.8 157.32 309.51 ;
   RECT 23.18 309.51 157.32 311.22 ;
   RECT 23.18 311.22 157.32 312.93 ;
   RECT 23.18 312.93 157.32 314.64 ;
   RECT 23.18 314.64 157.32 316.35 ;
   RECT 23.18 316.35 157.32 318.06 ;
   RECT 23.18 318.06 157.32 319.77 ;
   RECT 23.18 319.77 157.32 321.48 ;
   RECT 23.18 321.48 157.32 323.19 ;
   RECT 23.18 323.19 157.32 324.9 ;
   RECT 23.18 324.9 157.32 326.61 ;
   RECT 23.18 326.61 157.32 328.32 ;
   RECT 23.18 328.32 157.32 330.03 ;
   RECT 23.18 330.03 157.32 331.74 ;
   RECT 23.18 331.74 157.32 333.45 ;
   RECT 23.18 333.45 157.32 335.16 ;
   RECT 23.18 335.16 157.32 336.87 ;
   RECT 23.18 336.87 157.32 338.58 ;
   RECT 23.18 338.58 157.32 340.29 ;
   RECT 23.18 340.29 157.32 342.0 ;
   RECT 23.18 342.0 157.32 343.71 ;
   RECT 23.18 343.71 157.32 345.42 ;
   RECT 23.18 345.42 157.32 347.13 ;
   RECT 23.18 347.13 157.32 348.84 ;
   RECT 23.18 348.84 157.32 350.55 ;
   RECT 23.18 350.55 157.32 352.26 ;
   RECT 23.18 352.26 157.32 353.97 ;
   RECT 23.18 353.97 157.32 355.68 ;
   RECT 0.0 355.68 157.32 357.39 ;
   RECT 0.0 357.39 157.32 359.1 ;
   RECT 0.0 359.1 157.32 360.81 ;
   RECT 0.0 360.81 157.32 362.52 ;
   RECT 0.0 362.52 157.32 364.23 ;
   RECT 0.0 364.23 157.32 365.94 ;
   RECT 0.0 365.94 157.32 367.65 ;
   RECT 0.0 367.65 157.32 369.36 ;
   RECT 0.0 369.36 157.32 371.07 ;
   RECT 0.0 371.07 157.32 372.78 ;
   RECT 0.0 372.78 157.32 374.49 ;
   RECT 0.0 374.49 157.32 376.2 ;
   RECT 0.0 376.2 157.32 377.91 ;
   RECT 0.0 377.91 157.32 379.62 ;
   RECT 0.0 379.62 157.32 381.33 ;
   RECT 0.0 381.33 157.32 383.04 ;
   RECT 0.0 383.04 157.32 384.75 ;
   RECT 23.18 384.75 157.32 386.46 ;
   RECT 23.18 386.46 157.32 388.17 ;
   RECT 23.18 388.17 157.32 389.88 ;
   RECT 23.18 389.88 157.32 391.59 ;
   RECT 23.18 391.59 157.32 393.3 ;
   RECT 23.18 393.3 157.32 395.01 ;
   RECT 23.18 395.01 157.32 396.72 ;
   RECT 23.18 396.72 157.32 398.43 ;
   RECT 23.18 398.43 157.32 400.14 ;
   RECT 23.18 400.14 157.32 401.85 ;
   RECT 23.18 401.85 157.32 403.56 ;
   RECT 23.18 403.56 157.32 405.27 ;
   RECT 23.18 405.27 157.32 406.98 ;
   RECT 23.18 406.98 157.32 408.69 ;
   RECT 23.18 408.69 157.32 410.4 ;
   RECT 23.18 410.4 157.32 412.11 ;
   RECT 23.18 412.11 157.32 413.82 ;
   RECT 23.18 413.82 157.32 415.53 ;
   RECT 23.18 415.53 157.32 417.24 ;
   RECT 23.18 417.24 157.32 418.95 ;
   RECT 23.18 418.95 157.32 420.66 ;
   RECT 23.18 420.66 157.32 422.37 ;
   RECT 23.18 422.37 157.32 424.08 ;
   RECT 23.18 424.08 157.32 425.79 ;
   RECT 23.18 425.79 157.32 427.5 ;
   RECT 23.18 427.5 157.32 429.21 ;
   RECT 23.18 429.21 157.32 430.92 ;
   RECT 23.18 430.92 157.32 432.63 ;
   RECT 23.18 432.63 157.32 434.34 ;
   RECT 23.18 434.34 157.32 436.05 ;
   RECT 23.18 436.05 157.32 437.76 ;
   RECT 23.18 437.76 157.32 439.47 ;
   RECT 23.18 439.47 157.32 441.18 ;
   RECT 23.18 441.18 157.32 442.89 ;
   RECT 23.18 442.89 157.32 444.6 ;
   RECT 23.18 444.6 157.32 446.31 ;
   RECT 23.18 446.31 157.32 448.02 ;
   RECT 23.18 448.02 157.32 449.73 ;
   RECT 23.18 449.73 157.32 451.44 ;
   RECT 23.18 451.44 157.32 453.15 ;
   RECT 23.18 453.15 157.32 454.86 ;
   RECT 23.18 454.86 157.32 456.57 ;
   RECT 23.18 456.57 157.32 458.28 ;
   RECT 23.18 458.28 157.32 459.99 ;
   RECT 23.18 459.99 157.32 461.7 ;
   RECT 23.18 461.7 157.32 463.41 ;
   RECT 23.18 463.41 157.32 465.12 ;
   RECT 23.18 465.12 157.32 466.83 ;
   RECT 23.18 466.83 157.32 468.54 ;
   RECT 23.18 468.54 157.32 470.25 ;
   RECT 23.18 470.25 157.32 471.96 ;
   RECT 23.18 471.96 157.32 473.67 ;
   RECT 23.18 473.67 157.32 475.38 ;
   RECT 23.18 475.38 157.32 477.09 ;
   RECT 23.18 477.09 157.32 478.8 ;
   RECT 23.18 478.8 157.32 480.51 ;
   RECT 23.18 480.51 157.32 482.22 ;
   RECT 23.18 482.22 157.32 483.93 ;
   RECT 23.18 483.93 157.32 485.64 ;
   RECT 23.18 485.64 157.32 487.35 ;
   RECT 23.18 487.35 157.32 489.06 ;
   RECT 23.18 489.06 157.32 490.77 ;
   RECT 23.18 490.77 157.32 492.48 ;
   RECT 23.18 492.48 157.32 494.19 ;
   RECT 23.18 494.19 157.32 495.9 ;
   RECT 23.18 495.9 157.32 497.61 ;
   RECT 23.18 497.61 157.32 499.32 ;
   RECT 23.18 499.32 157.32 501.03 ;
   RECT 23.18 501.03 157.32 502.74 ;
   RECT 23.18 502.74 157.32 504.45 ;
   RECT 23.18 504.45 157.32 506.16 ;
   RECT 23.18 506.16 157.32 507.87 ;
   RECT 23.18 507.87 157.32 509.58 ;
   RECT 23.18 509.58 157.32 511.29 ;
   RECT 23.18 511.29 157.32 513.0 ;
   RECT 23.18 513.0 157.32 514.71 ;
   RECT 23.18 514.71 157.32 516.42 ;
   RECT 23.18 516.42 157.32 518.13 ;
   RECT 23.18 518.13 157.32 519.84 ;
   RECT 23.18 519.84 157.32 521.55 ;
   RECT 23.18 521.55 157.32 523.26 ;
   RECT 23.18 523.26 157.32 524.97 ;
   RECT 23.18 524.97 157.32 526.68 ;
   RECT 23.18 526.68 157.32 528.39 ;
   RECT 23.18 528.39 157.32 530.1 ;
   RECT 23.18 530.1 157.32 531.81 ;
   RECT 23.18 531.81 157.32 533.52 ;
   RECT 23.18 533.52 157.32 535.23 ;
   RECT 23.18 535.23 157.32 536.94 ;
   RECT 23.18 536.94 157.32 538.65 ;
   RECT 23.18 538.65 157.32 540.36 ;
   RECT 23.18 540.36 157.32 542.07 ;
   RECT 23.18 542.07 157.32 543.78 ;
   RECT 23.18 543.78 157.32 545.49 ;
   RECT 23.18 545.49 157.32 547.2 ;
   RECT 23.18 547.2 157.32 548.91 ;
   RECT 23.18 548.91 157.32 550.62 ;
   RECT 23.18 550.62 157.32 552.33 ;
   RECT 23.18 552.33 157.32 554.04 ;
   RECT 23.18 554.04 157.32 555.75 ;
   RECT 23.18 555.75 157.32 557.46 ;
   RECT 23.18 557.46 157.32 559.17 ;
   RECT 23.18 559.17 157.32 560.88 ;
   RECT 23.18 560.88 157.32 562.59 ;
   RECT 23.18 562.59 157.32 564.3 ;
   RECT 23.18 564.3 157.32 566.01 ;
   RECT 23.18 566.01 157.32 567.72 ;
   RECT 23.18 567.72 157.32 569.43 ;
   RECT 23.18 569.43 157.32 571.14 ;
   RECT 23.18 571.14 157.32 572.85 ;
   RECT 23.18 572.85 157.32 574.56 ;
   RECT 23.18 574.56 157.32 576.27 ;
   RECT 23.18 576.27 157.32 577.98 ;
   RECT 23.18 577.98 157.32 579.69 ;
   RECT 23.18 579.69 157.32 581.4 ;
   RECT 23.18 581.4 157.32 583.11 ;
   RECT 23.18 583.11 157.32 584.82 ;
   RECT 23.18 584.82 157.32 586.53 ;
   RECT 23.18 586.53 157.32 588.24 ;
   RECT 23.18 588.24 157.32 589.95 ;
   RECT 23.18 589.95 157.32 591.66 ;
   RECT 23.18 591.66 157.32 593.37 ;
   RECT 23.18 593.37 157.32 595.08 ;
   RECT 23.18 595.08 157.32 596.79 ;
   RECT 23.18 596.79 157.32 598.5 ;
   RECT 23.18 598.5 157.32 600.21 ;
   RECT 23.18 600.21 157.32 601.92 ;
   RECT 23.18 601.92 157.32 603.63 ;
   RECT 23.18 603.63 157.32 605.34 ;
   RECT 23.18 605.34 157.32 607.05 ;
   RECT 23.18 607.05 157.32 608.76 ;
   RECT 23.18 608.76 157.32 610.47 ;
   RECT 23.18 610.47 157.32 612.18 ;
   RECT 23.18 612.18 157.32 613.89 ;
   RECT 23.18 613.89 157.32 615.6 ;
   RECT 23.18 615.6 157.32 617.31 ;
   RECT 23.18 617.31 157.32 619.02 ;
   RECT 23.18 619.02 157.32 620.73 ;
   RECT 23.18 620.73 157.32 622.44 ;
   RECT 23.18 622.44 157.32 624.15 ;
   RECT 23.18 624.15 157.32 625.86 ;
   RECT 23.18 625.86 157.32 627.57 ;
   RECT 23.18 627.57 157.32 629.28 ;
   RECT 23.18 629.28 157.32 630.99 ;
   RECT 23.18 630.99 157.32 632.7 ;
   RECT 23.18 632.7 157.32 634.41 ;
   RECT 23.18 634.41 157.32 636.12 ;
   RECT 23.18 636.12 157.32 637.83 ;
   RECT 23.18 637.83 157.32 639.54 ;
   RECT 23.18 639.54 157.32 641.25 ;
   RECT 23.18 641.25 157.32 642.96 ;
   RECT 23.18 642.96 157.32 644.67 ;
   RECT 23.18 644.67 157.32 646.38 ;
   RECT 23.18 646.38 157.32 648.09 ;
   RECT 23.18 648.09 157.32 649.8 ;
   RECT 23.18 649.8 157.32 651.51 ;
   RECT 23.18 651.51 157.32 653.22 ;
   RECT 23.18 653.22 157.32 654.93 ;
   RECT 23.18 654.93 157.32 656.64 ;
   RECT 23.18 656.64 157.32 658.35 ;
   RECT 23.18 658.35 157.32 660.06 ;
   RECT 23.18 660.06 157.32 661.77 ;
   RECT 23.18 661.77 157.32 663.48 ;
   RECT 23.18 663.48 157.32 665.19 ;
   RECT 23.18 665.19 157.32 666.9 ;
   RECT 23.18 666.9 157.32 668.61 ;
   RECT 23.18 668.61 157.32 670.32 ;
   RECT 23.18 670.32 157.32 672.03 ;
   RECT 23.18 672.03 157.32 673.74 ;
   RECT 23.18 673.74 157.32 675.45 ;
   RECT 23.18 675.45 157.32 677.16 ;
   RECT 23.18 677.16 157.32 678.87 ;
   RECT 23.18 678.87 157.32 680.58 ;
   RECT 23.18 680.58 157.32 682.29 ;
   RECT 23.18 682.29 157.32 684.0 ;
   RECT 23.18 684.0 157.32 685.71 ;
   RECT 23.18 685.71 157.32 687.42 ;
   RECT 23.18 687.42 157.32 689.13 ;
   RECT 23.18 689.13 157.32 690.84 ;
   RECT 23.18 690.84 157.32 692.55 ;
   RECT 23.18 692.55 157.32 694.26 ;
   RECT 23.18 694.26 157.32 695.97 ;
   RECT 23.18 695.97 157.32 697.68 ;
   RECT 23.18 697.68 157.32 699.39 ;
   RECT 23.18 699.39 157.32 701.1 ;
   RECT 23.18 701.1 157.32 702.81 ;
   RECT 23.18 702.81 157.32 704.52 ;
   RECT 23.18 704.52 157.32 706.23 ;
   RECT 23.18 706.23 157.32 707.94 ;
   RECT 23.18 707.94 157.32 709.65 ;
   RECT 23.18 709.65 157.32 711.36 ;
   RECT 23.18 711.36 157.32 713.07 ;
   RECT 23.18 713.07 157.32 714.78 ;
   RECT 23.18 714.78 157.32 716.49 ;
   RECT 23.18 716.49 157.32 718.2 ;
   RECT 23.18 718.2 157.32 719.91 ;
   RECT 23.18 719.91 157.32 721.62 ;
   RECT 23.18 721.62 157.32 723.33 ;
   RECT 23.18 723.33 157.32 725.04 ;
   RECT 23.18 725.04 157.32 726.75 ;
   RECT 23.18 726.75 157.32 728.46 ;
   RECT 23.18 728.46 157.32 730.17 ;
   RECT 23.18 730.17 157.32 731.88 ;
   RECT 23.18 731.88 157.32 733.59 ;
   RECT 23.18 733.59 157.32 735.3 ;
   RECT 23.18 735.3 157.32 737.01 ;
   RECT 23.18 737.01 157.32 738.72 ;
   RECT 23.18 738.72 157.32 740.43 ;
   RECT 23.18 740.43 157.32 742.14 ;
   RECT 23.18 742.14 157.32 743.85 ;
   RECT 23.18 743.85 157.32 745.56 ;
   RECT 23.18 745.56 157.32 747.27 ;
   RECT 23.18 747.27 157.32 748.98 ;
   RECT 23.18 748.98 157.32 750.69 ;
   RECT 23.18 750.69 157.32 752.4 ;
   RECT 23.18 752.4 157.32 754.11 ;
  LAYER via2 ;
   RECT 23.18 0.0 157.32 1.71 ;
   RECT 23.18 1.71 157.32 3.42 ;
   RECT 23.18 3.42 157.32 5.13 ;
   RECT 23.18 5.13 157.32 6.84 ;
   RECT 23.18 6.84 157.32 8.55 ;
   RECT 23.18 8.55 157.32 10.26 ;
   RECT 23.18 10.26 157.32 11.97 ;
   RECT 23.18 11.97 157.32 13.68 ;
   RECT 23.18 13.68 157.32 15.39 ;
   RECT 23.18 15.39 157.32 17.1 ;
   RECT 23.18 17.1 157.32 18.81 ;
   RECT 23.18 18.81 157.32 20.52 ;
   RECT 23.18 20.52 157.32 22.23 ;
   RECT 23.18 22.23 157.32 23.94 ;
   RECT 23.18 23.94 157.32 25.65 ;
   RECT 23.18 25.65 157.32 27.36 ;
   RECT 23.18 27.36 157.32 29.07 ;
   RECT 23.18 29.07 157.32 30.78 ;
   RECT 23.18 30.78 157.32 32.49 ;
   RECT 23.18 32.49 157.32 34.2 ;
   RECT 23.18 34.2 157.32 35.91 ;
   RECT 23.18 35.91 157.32 37.62 ;
   RECT 23.18 37.62 157.32 39.33 ;
   RECT 23.18 39.33 157.32 41.04 ;
   RECT 23.18 41.04 157.32 42.75 ;
   RECT 23.18 42.75 157.32 44.46 ;
   RECT 23.18 44.46 157.32 46.17 ;
   RECT 23.18 46.17 157.32 47.88 ;
   RECT 23.18 47.88 157.32 49.59 ;
   RECT 23.18 49.59 157.32 51.3 ;
   RECT 23.18 51.3 157.32 53.01 ;
   RECT 23.18 53.01 157.32 54.72 ;
   RECT 23.18 54.72 157.32 56.43 ;
   RECT 23.18 56.43 157.32 58.14 ;
   RECT 23.18 58.14 157.32 59.85 ;
   RECT 23.18 59.85 157.32 61.56 ;
   RECT 23.18 61.56 157.32 63.27 ;
   RECT 23.18 63.27 157.32 64.98 ;
   RECT 23.18 64.98 157.32 66.69 ;
   RECT 23.18 66.69 157.32 68.4 ;
   RECT 23.18 68.4 157.32 70.11 ;
   RECT 23.18 70.11 157.32 71.82 ;
   RECT 23.18 71.82 157.32 73.53 ;
   RECT 23.18 73.53 157.32 75.24 ;
   RECT 23.18 75.24 157.32 76.95 ;
   RECT 23.18 76.95 157.32 78.66 ;
   RECT 23.18 78.66 157.32 80.37 ;
   RECT 23.18 80.37 157.32 82.08 ;
   RECT 23.18 82.08 157.32 83.79 ;
   RECT 23.18 83.79 157.32 85.5 ;
   RECT 23.18 85.5 157.32 87.21 ;
   RECT 23.18 87.21 157.32 88.92 ;
   RECT 23.18 88.92 157.32 90.63 ;
   RECT 23.18 90.63 157.32 92.34 ;
   RECT 23.18 92.34 157.32 94.05 ;
   RECT 23.18 94.05 157.32 95.76 ;
   RECT 23.18 95.76 157.32 97.47 ;
   RECT 23.18 97.47 157.32 99.18 ;
   RECT 23.18 99.18 157.32 100.89 ;
   RECT 23.18 100.89 157.32 102.6 ;
   RECT 23.18 102.6 157.32 104.31 ;
   RECT 23.18 104.31 157.32 106.02 ;
   RECT 23.18 106.02 157.32 107.73 ;
   RECT 23.18 107.73 157.32 109.44 ;
   RECT 23.18 109.44 157.32 111.15 ;
   RECT 23.18 111.15 157.32 112.86 ;
   RECT 23.18 112.86 157.32 114.57 ;
   RECT 23.18 114.57 157.32 116.28 ;
   RECT 23.18 116.28 157.32 117.99 ;
   RECT 23.18 117.99 157.32 119.7 ;
   RECT 23.18 119.7 157.32 121.41 ;
   RECT 23.18 121.41 157.32 123.12 ;
   RECT 23.18 123.12 157.32 124.83 ;
   RECT 23.18 124.83 157.32 126.54 ;
   RECT 23.18 126.54 157.32 128.25 ;
   RECT 23.18 128.25 157.32 129.96 ;
   RECT 23.18 129.96 157.32 131.67 ;
   RECT 23.18 131.67 157.32 133.38 ;
   RECT 23.18 133.38 157.32 135.09 ;
   RECT 23.18 135.09 157.32 136.8 ;
   RECT 23.18 136.8 157.32 138.51 ;
   RECT 23.18 138.51 157.32 140.22 ;
   RECT 23.18 140.22 157.32 141.93 ;
   RECT 23.18 141.93 157.32 143.64 ;
   RECT 23.18 143.64 157.32 145.35 ;
   RECT 23.18 145.35 157.32 147.06 ;
   RECT 23.18 147.06 157.32 148.77 ;
   RECT 23.18 148.77 157.32 150.48 ;
   RECT 23.18 150.48 157.32 152.19 ;
   RECT 23.18 152.19 157.32 153.9 ;
   RECT 23.18 153.9 157.32 155.61 ;
   RECT 23.18 155.61 157.32 157.32 ;
   RECT 23.18 157.32 157.32 159.03 ;
   RECT 23.18 159.03 157.32 160.74 ;
   RECT 23.18 160.74 157.32 162.45 ;
   RECT 23.18 162.45 157.32 164.16 ;
   RECT 23.18 164.16 157.32 165.87 ;
   RECT 23.18 165.87 157.32 167.58 ;
   RECT 23.18 167.58 157.32 169.29 ;
   RECT 23.18 169.29 157.32 171.0 ;
   RECT 23.18 171.0 157.32 172.71 ;
   RECT 23.18 172.71 157.32 174.42 ;
   RECT 23.18 174.42 157.32 176.13 ;
   RECT 23.18 176.13 157.32 177.84 ;
   RECT 23.18 177.84 157.32 179.55 ;
   RECT 23.18 179.55 157.32 181.26 ;
   RECT 23.18 181.26 157.32 182.97 ;
   RECT 23.18 182.97 157.32 184.68 ;
   RECT 23.18 184.68 157.32 186.39 ;
   RECT 23.18 186.39 157.32 188.1 ;
   RECT 23.18 188.1 157.32 189.81 ;
   RECT 23.18 189.81 157.32 191.52 ;
   RECT 23.18 191.52 157.32 193.23 ;
   RECT 23.18 193.23 157.32 194.94 ;
   RECT 23.18 194.94 157.32 196.65 ;
   RECT 23.18 196.65 157.32 198.36 ;
   RECT 23.18 198.36 157.32 200.07 ;
   RECT 23.18 200.07 157.32 201.78 ;
   RECT 23.18 201.78 157.32 203.49 ;
   RECT 23.18 203.49 157.32 205.2 ;
   RECT 23.18 205.2 157.32 206.91 ;
   RECT 23.18 206.91 157.32 208.62 ;
   RECT 23.18 208.62 157.32 210.33 ;
   RECT 23.18 210.33 157.32 212.04 ;
   RECT 23.18 212.04 157.32 213.75 ;
   RECT 23.18 213.75 157.32 215.46 ;
   RECT 23.18 215.46 157.32 217.17 ;
   RECT 23.18 217.17 157.32 218.88 ;
   RECT 23.18 218.88 157.32 220.59 ;
   RECT 23.18 220.59 157.32 222.3 ;
   RECT 23.18 222.3 157.32 224.01 ;
   RECT 23.18 224.01 157.32 225.72 ;
   RECT 23.18 225.72 157.32 227.43 ;
   RECT 23.18 227.43 157.32 229.14 ;
   RECT 23.18 229.14 157.32 230.85 ;
   RECT 23.18 230.85 157.32 232.56 ;
   RECT 23.18 232.56 157.32 234.27 ;
   RECT 23.18 234.27 157.32 235.98 ;
   RECT 23.18 235.98 157.32 237.69 ;
   RECT 23.18 237.69 157.32 239.4 ;
   RECT 23.18 239.4 157.32 241.11 ;
   RECT 23.18 241.11 157.32 242.82 ;
   RECT 23.18 242.82 157.32 244.53 ;
   RECT 23.18 244.53 157.32 246.24 ;
   RECT 23.18 246.24 157.32 247.95 ;
   RECT 23.18 247.95 157.32 249.66 ;
   RECT 23.18 249.66 157.32 251.37 ;
   RECT 23.18 251.37 157.32 253.08 ;
   RECT 23.18 253.08 157.32 254.79 ;
   RECT 23.18 254.79 157.32 256.5 ;
   RECT 23.18 256.5 157.32 258.21 ;
   RECT 23.18 258.21 157.32 259.92 ;
   RECT 23.18 259.92 157.32 261.63 ;
   RECT 23.18 261.63 157.32 263.34 ;
   RECT 23.18 263.34 157.32 265.05 ;
   RECT 23.18 265.05 157.32 266.76 ;
   RECT 23.18 266.76 157.32 268.47 ;
   RECT 23.18 268.47 157.32 270.18 ;
   RECT 23.18 270.18 157.32 271.89 ;
   RECT 23.18 271.89 157.32 273.6 ;
   RECT 23.18 273.6 157.32 275.31 ;
   RECT 23.18 275.31 157.32 277.02 ;
   RECT 23.18 277.02 157.32 278.73 ;
   RECT 23.18 278.73 157.32 280.44 ;
   RECT 23.18 280.44 157.32 282.15 ;
   RECT 23.18 282.15 157.32 283.86 ;
   RECT 23.18 283.86 157.32 285.57 ;
   RECT 23.18 285.57 157.32 287.28 ;
   RECT 23.18 287.28 157.32 288.99 ;
   RECT 23.18 288.99 157.32 290.7 ;
   RECT 23.18 290.7 157.32 292.41 ;
   RECT 23.18 292.41 157.32 294.12 ;
   RECT 23.18 294.12 157.32 295.83 ;
   RECT 23.18 295.83 157.32 297.54 ;
   RECT 23.18 297.54 157.32 299.25 ;
   RECT 23.18 299.25 157.32 300.96 ;
   RECT 23.18 300.96 157.32 302.67 ;
   RECT 23.18 302.67 157.32 304.38 ;
   RECT 23.18 304.38 157.32 306.09 ;
   RECT 23.18 306.09 157.32 307.8 ;
   RECT 23.18 307.8 157.32 309.51 ;
   RECT 23.18 309.51 157.32 311.22 ;
   RECT 23.18 311.22 157.32 312.93 ;
   RECT 23.18 312.93 157.32 314.64 ;
   RECT 23.18 314.64 157.32 316.35 ;
   RECT 23.18 316.35 157.32 318.06 ;
   RECT 23.18 318.06 157.32 319.77 ;
   RECT 23.18 319.77 157.32 321.48 ;
   RECT 23.18 321.48 157.32 323.19 ;
   RECT 23.18 323.19 157.32 324.9 ;
   RECT 23.18 324.9 157.32 326.61 ;
   RECT 23.18 326.61 157.32 328.32 ;
   RECT 23.18 328.32 157.32 330.03 ;
   RECT 23.18 330.03 157.32 331.74 ;
   RECT 23.18 331.74 157.32 333.45 ;
   RECT 23.18 333.45 157.32 335.16 ;
   RECT 23.18 335.16 157.32 336.87 ;
   RECT 23.18 336.87 157.32 338.58 ;
   RECT 23.18 338.58 157.32 340.29 ;
   RECT 23.18 340.29 157.32 342.0 ;
   RECT 23.18 342.0 157.32 343.71 ;
   RECT 23.18 343.71 157.32 345.42 ;
   RECT 23.18 345.42 157.32 347.13 ;
   RECT 23.18 347.13 157.32 348.84 ;
   RECT 23.18 348.84 157.32 350.55 ;
   RECT 23.18 350.55 157.32 352.26 ;
   RECT 23.18 352.26 157.32 353.97 ;
   RECT 23.18 353.97 157.32 355.68 ;
   RECT 0.0 355.68 157.32 357.39 ;
   RECT 0.0 357.39 157.32 359.1 ;
   RECT 0.0 359.1 157.32 360.81 ;
   RECT 0.0 360.81 157.32 362.52 ;
   RECT 0.0 362.52 157.32 364.23 ;
   RECT 0.0 364.23 157.32 365.94 ;
   RECT 0.0 365.94 157.32 367.65 ;
   RECT 0.0 367.65 157.32 369.36 ;
   RECT 0.0 369.36 157.32 371.07 ;
   RECT 0.0 371.07 157.32 372.78 ;
   RECT 0.0 372.78 157.32 374.49 ;
   RECT 0.0 374.49 157.32 376.2 ;
   RECT 0.0 376.2 157.32 377.91 ;
   RECT 0.0 377.91 157.32 379.62 ;
   RECT 0.0 379.62 157.32 381.33 ;
   RECT 0.0 381.33 157.32 383.04 ;
   RECT 0.0 383.04 157.32 384.75 ;
   RECT 23.18 384.75 157.32 386.46 ;
   RECT 23.18 386.46 157.32 388.17 ;
   RECT 23.18 388.17 157.32 389.88 ;
   RECT 23.18 389.88 157.32 391.59 ;
   RECT 23.18 391.59 157.32 393.3 ;
   RECT 23.18 393.3 157.32 395.01 ;
   RECT 23.18 395.01 157.32 396.72 ;
   RECT 23.18 396.72 157.32 398.43 ;
   RECT 23.18 398.43 157.32 400.14 ;
   RECT 23.18 400.14 157.32 401.85 ;
   RECT 23.18 401.85 157.32 403.56 ;
   RECT 23.18 403.56 157.32 405.27 ;
   RECT 23.18 405.27 157.32 406.98 ;
   RECT 23.18 406.98 157.32 408.69 ;
   RECT 23.18 408.69 157.32 410.4 ;
   RECT 23.18 410.4 157.32 412.11 ;
   RECT 23.18 412.11 157.32 413.82 ;
   RECT 23.18 413.82 157.32 415.53 ;
   RECT 23.18 415.53 157.32 417.24 ;
   RECT 23.18 417.24 157.32 418.95 ;
   RECT 23.18 418.95 157.32 420.66 ;
   RECT 23.18 420.66 157.32 422.37 ;
   RECT 23.18 422.37 157.32 424.08 ;
   RECT 23.18 424.08 157.32 425.79 ;
   RECT 23.18 425.79 157.32 427.5 ;
   RECT 23.18 427.5 157.32 429.21 ;
   RECT 23.18 429.21 157.32 430.92 ;
   RECT 23.18 430.92 157.32 432.63 ;
   RECT 23.18 432.63 157.32 434.34 ;
   RECT 23.18 434.34 157.32 436.05 ;
   RECT 23.18 436.05 157.32 437.76 ;
   RECT 23.18 437.76 157.32 439.47 ;
   RECT 23.18 439.47 157.32 441.18 ;
   RECT 23.18 441.18 157.32 442.89 ;
   RECT 23.18 442.89 157.32 444.6 ;
   RECT 23.18 444.6 157.32 446.31 ;
   RECT 23.18 446.31 157.32 448.02 ;
   RECT 23.18 448.02 157.32 449.73 ;
   RECT 23.18 449.73 157.32 451.44 ;
   RECT 23.18 451.44 157.32 453.15 ;
   RECT 23.18 453.15 157.32 454.86 ;
   RECT 23.18 454.86 157.32 456.57 ;
   RECT 23.18 456.57 157.32 458.28 ;
   RECT 23.18 458.28 157.32 459.99 ;
   RECT 23.18 459.99 157.32 461.7 ;
   RECT 23.18 461.7 157.32 463.41 ;
   RECT 23.18 463.41 157.32 465.12 ;
   RECT 23.18 465.12 157.32 466.83 ;
   RECT 23.18 466.83 157.32 468.54 ;
   RECT 23.18 468.54 157.32 470.25 ;
   RECT 23.18 470.25 157.32 471.96 ;
   RECT 23.18 471.96 157.32 473.67 ;
   RECT 23.18 473.67 157.32 475.38 ;
   RECT 23.18 475.38 157.32 477.09 ;
   RECT 23.18 477.09 157.32 478.8 ;
   RECT 23.18 478.8 157.32 480.51 ;
   RECT 23.18 480.51 157.32 482.22 ;
   RECT 23.18 482.22 157.32 483.93 ;
   RECT 23.18 483.93 157.32 485.64 ;
   RECT 23.18 485.64 157.32 487.35 ;
   RECT 23.18 487.35 157.32 489.06 ;
   RECT 23.18 489.06 157.32 490.77 ;
   RECT 23.18 490.77 157.32 492.48 ;
   RECT 23.18 492.48 157.32 494.19 ;
   RECT 23.18 494.19 157.32 495.9 ;
   RECT 23.18 495.9 157.32 497.61 ;
   RECT 23.18 497.61 157.32 499.32 ;
   RECT 23.18 499.32 157.32 501.03 ;
   RECT 23.18 501.03 157.32 502.74 ;
   RECT 23.18 502.74 157.32 504.45 ;
   RECT 23.18 504.45 157.32 506.16 ;
   RECT 23.18 506.16 157.32 507.87 ;
   RECT 23.18 507.87 157.32 509.58 ;
   RECT 23.18 509.58 157.32 511.29 ;
   RECT 23.18 511.29 157.32 513.0 ;
   RECT 23.18 513.0 157.32 514.71 ;
   RECT 23.18 514.71 157.32 516.42 ;
   RECT 23.18 516.42 157.32 518.13 ;
   RECT 23.18 518.13 157.32 519.84 ;
   RECT 23.18 519.84 157.32 521.55 ;
   RECT 23.18 521.55 157.32 523.26 ;
   RECT 23.18 523.26 157.32 524.97 ;
   RECT 23.18 524.97 157.32 526.68 ;
   RECT 23.18 526.68 157.32 528.39 ;
   RECT 23.18 528.39 157.32 530.1 ;
   RECT 23.18 530.1 157.32 531.81 ;
   RECT 23.18 531.81 157.32 533.52 ;
   RECT 23.18 533.52 157.32 535.23 ;
   RECT 23.18 535.23 157.32 536.94 ;
   RECT 23.18 536.94 157.32 538.65 ;
   RECT 23.18 538.65 157.32 540.36 ;
   RECT 23.18 540.36 157.32 542.07 ;
   RECT 23.18 542.07 157.32 543.78 ;
   RECT 23.18 543.78 157.32 545.49 ;
   RECT 23.18 545.49 157.32 547.2 ;
   RECT 23.18 547.2 157.32 548.91 ;
   RECT 23.18 548.91 157.32 550.62 ;
   RECT 23.18 550.62 157.32 552.33 ;
   RECT 23.18 552.33 157.32 554.04 ;
   RECT 23.18 554.04 157.32 555.75 ;
   RECT 23.18 555.75 157.32 557.46 ;
   RECT 23.18 557.46 157.32 559.17 ;
   RECT 23.18 559.17 157.32 560.88 ;
   RECT 23.18 560.88 157.32 562.59 ;
   RECT 23.18 562.59 157.32 564.3 ;
   RECT 23.18 564.3 157.32 566.01 ;
   RECT 23.18 566.01 157.32 567.72 ;
   RECT 23.18 567.72 157.32 569.43 ;
   RECT 23.18 569.43 157.32 571.14 ;
   RECT 23.18 571.14 157.32 572.85 ;
   RECT 23.18 572.85 157.32 574.56 ;
   RECT 23.18 574.56 157.32 576.27 ;
   RECT 23.18 576.27 157.32 577.98 ;
   RECT 23.18 577.98 157.32 579.69 ;
   RECT 23.18 579.69 157.32 581.4 ;
   RECT 23.18 581.4 157.32 583.11 ;
   RECT 23.18 583.11 157.32 584.82 ;
   RECT 23.18 584.82 157.32 586.53 ;
   RECT 23.18 586.53 157.32 588.24 ;
   RECT 23.18 588.24 157.32 589.95 ;
   RECT 23.18 589.95 157.32 591.66 ;
   RECT 23.18 591.66 157.32 593.37 ;
   RECT 23.18 593.37 157.32 595.08 ;
   RECT 23.18 595.08 157.32 596.79 ;
   RECT 23.18 596.79 157.32 598.5 ;
   RECT 23.18 598.5 157.32 600.21 ;
   RECT 23.18 600.21 157.32 601.92 ;
   RECT 23.18 601.92 157.32 603.63 ;
   RECT 23.18 603.63 157.32 605.34 ;
   RECT 23.18 605.34 157.32 607.05 ;
   RECT 23.18 607.05 157.32 608.76 ;
   RECT 23.18 608.76 157.32 610.47 ;
   RECT 23.18 610.47 157.32 612.18 ;
   RECT 23.18 612.18 157.32 613.89 ;
   RECT 23.18 613.89 157.32 615.6 ;
   RECT 23.18 615.6 157.32 617.31 ;
   RECT 23.18 617.31 157.32 619.02 ;
   RECT 23.18 619.02 157.32 620.73 ;
   RECT 23.18 620.73 157.32 622.44 ;
   RECT 23.18 622.44 157.32 624.15 ;
   RECT 23.18 624.15 157.32 625.86 ;
   RECT 23.18 625.86 157.32 627.57 ;
   RECT 23.18 627.57 157.32 629.28 ;
   RECT 23.18 629.28 157.32 630.99 ;
   RECT 23.18 630.99 157.32 632.7 ;
   RECT 23.18 632.7 157.32 634.41 ;
   RECT 23.18 634.41 157.32 636.12 ;
   RECT 23.18 636.12 157.32 637.83 ;
   RECT 23.18 637.83 157.32 639.54 ;
   RECT 23.18 639.54 157.32 641.25 ;
   RECT 23.18 641.25 157.32 642.96 ;
   RECT 23.18 642.96 157.32 644.67 ;
   RECT 23.18 644.67 157.32 646.38 ;
   RECT 23.18 646.38 157.32 648.09 ;
   RECT 23.18 648.09 157.32 649.8 ;
   RECT 23.18 649.8 157.32 651.51 ;
   RECT 23.18 651.51 157.32 653.22 ;
   RECT 23.18 653.22 157.32 654.93 ;
   RECT 23.18 654.93 157.32 656.64 ;
   RECT 23.18 656.64 157.32 658.35 ;
   RECT 23.18 658.35 157.32 660.06 ;
   RECT 23.18 660.06 157.32 661.77 ;
   RECT 23.18 661.77 157.32 663.48 ;
   RECT 23.18 663.48 157.32 665.19 ;
   RECT 23.18 665.19 157.32 666.9 ;
   RECT 23.18 666.9 157.32 668.61 ;
   RECT 23.18 668.61 157.32 670.32 ;
   RECT 23.18 670.32 157.32 672.03 ;
   RECT 23.18 672.03 157.32 673.74 ;
   RECT 23.18 673.74 157.32 675.45 ;
   RECT 23.18 675.45 157.32 677.16 ;
   RECT 23.18 677.16 157.32 678.87 ;
   RECT 23.18 678.87 157.32 680.58 ;
   RECT 23.18 680.58 157.32 682.29 ;
   RECT 23.18 682.29 157.32 684.0 ;
   RECT 23.18 684.0 157.32 685.71 ;
   RECT 23.18 685.71 157.32 687.42 ;
   RECT 23.18 687.42 157.32 689.13 ;
   RECT 23.18 689.13 157.32 690.84 ;
   RECT 23.18 690.84 157.32 692.55 ;
   RECT 23.18 692.55 157.32 694.26 ;
   RECT 23.18 694.26 157.32 695.97 ;
   RECT 23.18 695.97 157.32 697.68 ;
   RECT 23.18 697.68 157.32 699.39 ;
   RECT 23.18 699.39 157.32 701.1 ;
   RECT 23.18 701.1 157.32 702.81 ;
   RECT 23.18 702.81 157.32 704.52 ;
   RECT 23.18 704.52 157.32 706.23 ;
   RECT 23.18 706.23 157.32 707.94 ;
   RECT 23.18 707.94 157.32 709.65 ;
   RECT 23.18 709.65 157.32 711.36 ;
   RECT 23.18 711.36 157.32 713.07 ;
   RECT 23.18 713.07 157.32 714.78 ;
   RECT 23.18 714.78 157.32 716.49 ;
   RECT 23.18 716.49 157.32 718.2 ;
   RECT 23.18 718.2 157.32 719.91 ;
   RECT 23.18 719.91 157.32 721.62 ;
   RECT 23.18 721.62 157.32 723.33 ;
   RECT 23.18 723.33 157.32 725.04 ;
   RECT 23.18 725.04 157.32 726.75 ;
   RECT 23.18 726.75 157.32 728.46 ;
   RECT 23.18 728.46 157.32 730.17 ;
   RECT 23.18 730.17 157.32 731.88 ;
   RECT 23.18 731.88 157.32 733.59 ;
   RECT 23.18 733.59 157.32 735.3 ;
   RECT 23.18 735.3 157.32 737.01 ;
   RECT 23.18 737.01 157.32 738.72 ;
   RECT 23.18 738.72 157.32 740.43 ;
   RECT 23.18 740.43 157.32 742.14 ;
   RECT 23.18 742.14 157.32 743.85 ;
   RECT 23.18 743.85 157.32 745.56 ;
   RECT 23.18 745.56 157.32 747.27 ;
   RECT 23.18 747.27 157.32 748.98 ;
   RECT 23.18 748.98 157.32 750.69 ;
   RECT 23.18 750.69 157.32 752.4 ;
   RECT 23.18 752.4 157.32 754.11 ;
  LAYER metal3 ;
   RECT 23.18 0.0 157.32 1.71 ;
   RECT 23.18 1.71 157.32 3.42 ;
   RECT 23.18 3.42 157.32 5.13 ;
   RECT 23.18 5.13 157.32 6.84 ;
   RECT 23.18 6.84 157.32 8.55 ;
   RECT 23.18 8.55 157.32 10.26 ;
   RECT 23.18 10.26 157.32 11.97 ;
   RECT 23.18 11.97 157.32 13.68 ;
   RECT 23.18 13.68 157.32 15.39 ;
   RECT 23.18 15.39 157.32 17.1 ;
   RECT 23.18 17.1 157.32 18.81 ;
   RECT 23.18 18.81 157.32 20.52 ;
   RECT 23.18 20.52 157.32 22.23 ;
   RECT 23.18 22.23 157.32 23.94 ;
   RECT 23.18 23.94 157.32 25.65 ;
   RECT 23.18 25.65 157.32 27.36 ;
   RECT 23.18 27.36 157.32 29.07 ;
   RECT 23.18 29.07 157.32 30.78 ;
   RECT 23.18 30.78 157.32 32.49 ;
   RECT 23.18 32.49 157.32 34.2 ;
   RECT 23.18 34.2 157.32 35.91 ;
   RECT 23.18 35.91 157.32 37.62 ;
   RECT 23.18 37.62 157.32 39.33 ;
   RECT 23.18 39.33 157.32 41.04 ;
   RECT 23.18 41.04 157.32 42.75 ;
   RECT 23.18 42.75 157.32 44.46 ;
   RECT 23.18 44.46 157.32 46.17 ;
   RECT 23.18 46.17 157.32 47.88 ;
   RECT 23.18 47.88 157.32 49.59 ;
   RECT 23.18 49.59 157.32 51.3 ;
   RECT 23.18 51.3 157.32 53.01 ;
   RECT 23.18 53.01 157.32 54.72 ;
   RECT 23.18 54.72 157.32 56.43 ;
   RECT 23.18 56.43 157.32 58.14 ;
   RECT 23.18 58.14 157.32 59.85 ;
   RECT 23.18 59.85 157.32 61.56 ;
   RECT 23.18 61.56 157.32 63.27 ;
   RECT 23.18 63.27 157.32 64.98 ;
   RECT 23.18 64.98 157.32 66.69 ;
   RECT 23.18 66.69 157.32 68.4 ;
   RECT 23.18 68.4 157.32 70.11 ;
   RECT 23.18 70.11 157.32 71.82 ;
   RECT 23.18 71.82 157.32 73.53 ;
   RECT 23.18 73.53 157.32 75.24 ;
   RECT 23.18 75.24 157.32 76.95 ;
   RECT 23.18 76.95 157.32 78.66 ;
   RECT 23.18 78.66 157.32 80.37 ;
   RECT 23.18 80.37 157.32 82.08 ;
   RECT 23.18 82.08 157.32 83.79 ;
   RECT 23.18 83.79 157.32 85.5 ;
   RECT 23.18 85.5 157.32 87.21 ;
   RECT 23.18 87.21 157.32 88.92 ;
   RECT 23.18 88.92 157.32 90.63 ;
   RECT 23.18 90.63 157.32 92.34 ;
   RECT 23.18 92.34 157.32 94.05 ;
   RECT 23.18 94.05 157.32 95.76 ;
   RECT 23.18 95.76 157.32 97.47 ;
   RECT 23.18 97.47 157.32 99.18 ;
   RECT 23.18 99.18 157.32 100.89 ;
   RECT 23.18 100.89 157.32 102.6 ;
   RECT 23.18 102.6 157.32 104.31 ;
   RECT 23.18 104.31 157.32 106.02 ;
   RECT 23.18 106.02 157.32 107.73 ;
   RECT 23.18 107.73 157.32 109.44 ;
   RECT 23.18 109.44 157.32 111.15 ;
   RECT 23.18 111.15 157.32 112.86 ;
   RECT 23.18 112.86 157.32 114.57 ;
   RECT 23.18 114.57 157.32 116.28 ;
   RECT 23.18 116.28 157.32 117.99 ;
   RECT 23.18 117.99 157.32 119.7 ;
   RECT 23.18 119.7 157.32 121.41 ;
   RECT 23.18 121.41 157.32 123.12 ;
   RECT 23.18 123.12 157.32 124.83 ;
   RECT 23.18 124.83 157.32 126.54 ;
   RECT 23.18 126.54 157.32 128.25 ;
   RECT 23.18 128.25 157.32 129.96 ;
   RECT 23.18 129.96 157.32 131.67 ;
   RECT 23.18 131.67 157.32 133.38 ;
   RECT 23.18 133.38 157.32 135.09 ;
   RECT 23.18 135.09 157.32 136.8 ;
   RECT 23.18 136.8 157.32 138.51 ;
   RECT 23.18 138.51 157.32 140.22 ;
   RECT 23.18 140.22 157.32 141.93 ;
   RECT 23.18 141.93 157.32 143.64 ;
   RECT 23.18 143.64 157.32 145.35 ;
   RECT 23.18 145.35 157.32 147.06 ;
   RECT 23.18 147.06 157.32 148.77 ;
   RECT 23.18 148.77 157.32 150.48 ;
   RECT 23.18 150.48 157.32 152.19 ;
   RECT 23.18 152.19 157.32 153.9 ;
   RECT 23.18 153.9 157.32 155.61 ;
   RECT 23.18 155.61 157.32 157.32 ;
   RECT 23.18 157.32 157.32 159.03 ;
   RECT 23.18 159.03 157.32 160.74 ;
   RECT 23.18 160.74 157.32 162.45 ;
   RECT 23.18 162.45 157.32 164.16 ;
   RECT 23.18 164.16 157.32 165.87 ;
   RECT 23.18 165.87 157.32 167.58 ;
   RECT 23.18 167.58 157.32 169.29 ;
   RECT 23.18 169.29 157.32 171.0 ;
   RECT 23.18 171.0 157.32 172.71 ;
   RECT 23.18 172.71 157.32 174.42 ;
   RECT 23.18 174.42 157.32 176.13 ;
   RECT 23.18 176.13 157.32 177.84 ;
   RECT 23.18 177.84 157.32 179.55 ;
   RECT 23.18 179.55 157.32 181.26 ;
   RECT 23.18 181.26 157.32 182.97 ;
   RECT 23.18 182.97 157.32 184.68 ;
   RECT 23.18 184.68 157.32 186.39 ;
   RECT 23.18 186.39 157.32 188.1 ;
   RECT 23.18 188.1 157.32 189.81 ;
   RECT 23.18 189.81 157.32 191.52 ;
   RECT 23.18 191.52 157.32 193.23 ;
   RECT 23.18 193.23 157.32 194.94 ;
   RECT 23.18 194.94 157.32 196.65 ;
   RECT 23.18 196.65 157.32 198.36 ;
   RECT 23.18 198.36 157.32 200.07 ;
   RECT 23.18 200.07 157.32 201.78 ;
   RECT 23.18 201.78 157.32 203.49 ;
   RECT 23.18 203.49 157.32 205.2 ;
   RECT 23.18 205.2 157.32 206.91 ;
   RECT 23.18 206.91 157.32 208.62 ;
   RECT 23.18 208.62 157.32 210.33 ;
   RECT 23.18 210.33 157.32 212.04 ;
   RECT 23.18 212.04 157.32 213.75 ;
   RECT 23.18 213.75 157.32 215.46 ;
   RECT 23.18 215.46 157.32 217.17 ;
   RECT 23.18 217.17 157.32 218.88 ;
   RECT 23.18 218.88 157.32 220.59 ;
   RECT 23.18 220.59 157.32 222.3 ;
   RECT 23.18 222.3 157.32 224.01 ;
   RECT 23.18 224.01 157.32 225.72 ;
   RECT 23.18 225.72 157.32 227.43 ;
   RECT 23.18 227.43 157.32 229.14 ;
   RECT 23.18 229.14 157.32 230.85 ;
   RECT 23.18 230.85 157.32 232.56 ;
   RECT 23.18 232.56 157.32 234.27 ;
   RECT 23.18 234.27 157.32 235.98 ;
   RECT 23.18 235.98 157.32 237.69 ;
   RECT 23.18 237.69 157.32 239.4 ;
   RECT 23.18 239.4 157.32 241.11 ;
   RECT 23.18 241.11 157.32 242.82 ;
   RECT 23.18 242.82 157.32 244.53 ;
   RECT 23.18 244.53 157.32 246.24 ;
   RECT 23.18 246.24 157.32 247.95 ;
   RECT 23.18 247.95 157.32 249.66 ;
   RECT 23.18 249.66 157.32 251.37 ;
   RECT 23.18 251.37 157.32 253.08 ;
   RECT 23.18 253.08 157.32 254.79 ;
   RECT 23.18 254.79 157.32 256.5 ;
   RECT 23.18 256.5 157.32 258.21 ;
   RECT 23.18 258.21 157.32 259.92 ;
   RECT 23.18 259.92 157.32 261.63 ;
   RECT 23.18 261.63 157.32 263.34 ;
   RECT 23.18 263.34 157.32 265.05 ;
   RECT 23.18 265.05 157.32 266.76 ;
   RECT 23.18 266.76 157.32 268.47 ;
   RECT 23.18 268.47 157.32 270.18 ;
   RECT 23.18 270.18 157.32 271.89 ;
   RECT 23.18 271.89 157.32 273.6 ;
   RECT 23.18 273.6 157.32 275.31 ;
   RECT 23.18 275.31 157.32 277.02 ;
   RECT 23.18 277.02 157.32 278.73 ;
   RECT 23.18 278.73 157.32 280.44 ;
   RECT 23.18 280.44 157.32 282.15 ;
   RECT 23.18 282.15 157.32 283.86 ;
   RECT 23.18 283.86 157.32 285.57 ;
   RECT 23.18 285.57 157.32 287.28 ;
   RECT 23.18 287.28 157.32 288.99 ;
   RECT 23.18 288.99 157.32 290.7 ;
   RECT 23.18 290.7 157.32 292.41 ;
   RECT 23.18 292.41 157.32 294.12 ;
   RECT 23.18 294.12 157.32 295.83 ;
   RECT 23.18 295.83 157.32 297.54 ;
   RECT 23.18 297.54 157.32 299.25 ;
   RECT 23.18 299.25 157.32 300.96 ;
   RECT 23.18 300.96 157.32 302.67 ;
   RECT 23.18 302.67 157.32 304.38 ;
   RECT 23.18 304.38 157.32 306.09 ;
   RECT 23.18 306.09 157.32 307.8 ;
   RECT 23.18 307.8 157.32 309.51 ;
   RECT 23.18 309.51 157.32 311.22 ;
   RECT 23.18 311.22 157.32 312.93 ;
   RECT 23.18 312.93 157.32 314.64 ;
   RECT 23.18 314.64 157.32 316.35 ;
   RECT 23.18 316.35 157.32 318.06 ;
   RECT 23.18 318.06 157.32 319.77 ;
   RECT 23.18 319.77 157.32 321.48 ;
   RECT 23.18 321.48 157.32 323.19 ;
   RECT 23.18 323.19 157.32 324.9 ;
   RECT 23.18 324.9 157.32 326.61 ;
   RECT 23.18 326.61 157.32 328.32 ;
   RECT 23.18 328.32 157.32 330.03 ;
   RECT 23.18 330.03 157.32 331.74 ;
   RECT 23.18 331.74 157.32 333.45 ;
   RECT 23.18 333.45 157.32 335.16 ;
   RECT 23.18 335.16 157.32 336.87 ;
   RECT 23.18 336.87 157.32 338.58 ;
   RECT 23.18 338.58 157.32 340.29 ;
   RECT 23.18 340.29 157.32 342.0 ;
   RECT 23.18 342.0 157.32 343.71 ;
   RECT 23.18 343.71 157.32 345.42 ;
   RECT 23.18 345.42 157.32 347.13 ;
   RECT 23.18 347.13 157.32 348.84 ;
   RECT 23.18 348.84 157.32 350.55 ;
   RECT 23.18 350.55 157.32 352.26 ;
   RECT 23.18 352.26 157.32 353.97 ;
   RECT 23.18 353.97 157.32 355.68 ;
   RECT 0.0 355.68 157.32 357.39 ;
   RECT 0.0 357.39 157.32 359.1 ;
   RECT 0.0 359.1 157.32 360.81 ;
   RECT 0.0 360.81 157.32 362.52 ;
   RECT 0.0 362.52 157.32 364.23 ;
   RECT 0.0 364.23 157.32 365.94 ;
   RECT 0.0 365.94 157.32 367.65 ;
   RECT 0.0 367.65 157.32 369.36 ;
   RECT 0.0 369.36 157.32 371.07 ;
   RECT 0.0 371.07 157.32 372.78 ;
   RECT 0.0 372.78 157.32 374.49 ;
   RECT 0.0 374.49 157.32 376.2 ;
   RECT 0.0 376.2 157.32 377.91 ;
   RECT 0.0 377.91 157.32 379.62 ;
   RECT 0.0 379.62 157.32 381.33 ;
   RECT 0.0 381.33 157.32 383.04 ;
   RECT 0.0 383.04 157.32 384.75 ;
   RECT 23.18 384.75 157.32 386.46 ;
   RECT 23.18 386.46 157.32 388.17 ;
   RECT 23.18 388.17 157.32 389.88 ;
   RECT 23.18 389.88 157.32 391.59 ;
   RECT 23.18 391.59 157.32 393.3 ;
   RECT 23.18 393.3 157.32 395.01 ;
   RECT 23.18 395.01 157.32 396.72 ;
   RECT 23.18 396.72 157.32 398.43 ;
   RECT 23.18 398.43 157.32 400.14 ;
   RECT 23.18 400.14 157.32 401.85 ;
   RECT 23.18 401.85 157.32 403.56 ;
   RECT 23.18 403.56 157.32 405.27 ;
   RECT 23.18 405.27 157.32 406.98 ;
   RECT 23.18 406.98 157.32 408.69 ;
   RECT 23.18 408.69 157.32 410.4 ;
   RECT 23.18 410.4 157.32 412.11 ;
   RECT 23.18 412.11 157.32 413.82 ;
   RECT 23.18 413.82 157.32 415.53 ;
   RECT 23.18 415.53 157.32 417.24 ;
   RECT 23.18 417.24 157.32 418.95 ;
   RECT 23.18 418.95 157.32 420.66 ;
   RECT 23.18 420.66 157.32 422.37 ;
   RECT 23.18 422.37 157.32 424.08 ;
   RECT 23.18 424.08 157.32 425.79 ;
   RECT 23.18 425.79 157.32 427.5 ;
   RECT 23.18 427.5 157.32 429.21 ;
   RECT 23.18 429.21 157.32 430.92 ;
   RECT 23.18 430.92 157.32 432.63 ;
   RECT 23.18 432.63 157.32 434.34 ;
   RECT 23.18 434.34 157.32 436.05 ;
   RECT 23.18 436.05 157.32 437.76 ;
   RECT 23.18 437.76 157.32 439.47 ;
   RECT 23.18 439.47 157.32 441.18 ;
   RECT 23.18 441.18 157.32 442.89 ;
   RECT 23.18 442.89 157.32 444.6 ;
   RECT 23.18 444.6 157.32 446.31 ;
   RECT 23.18 446.31 157.32 448.02 ;
   RECT 23.18 448.02 157.32 449.73 ;
   RECT 23.18 449.73 157.32 451.44 ;
   RECT 23.18 451.44 157.32 453.15 ;
   RECT 23.18 453.15 157.32 454.86 ;
   RECT 23.18 454.86 157.32 456.57 ;
   RECT 23.18 456.57 157.32 458.28 ;
   RECT 23.18 458.28 157.32 459.99 ;
   RECT 23.18 459.99 157.32 461.7 ;
   RECT 23.18 461.7 157.32 463.41 ;
   RECT 23.18 463.41 157.32 465.12 ;
   RECT 23.18 465.12 157.32 466.83 ;
   RECT 23.18 466.83 157.32 468.54 ;
   RECT 23.18 468.54 157.32 470.25 ;
   RECT 23.18 470.25 157.32 471.96 ;
   RECT 23.18 471.96 157.32 473.67 ;
   RECT 23.18 473.67 157.32 475.38 ;
   RECT 23.18 475.38 157.32 477.09 ;
   RECT 23.18 477.09 157.32 478.8 ;
   RECT 23.18 478.8 157.32 480.51 ;
   RECT 23.18 480.51 157.32 482.22 ;
   RECT 23.18 482.22 157.32 483.93 ;
   RECT 23.18 483.93 157.32 485.64 ;
   RECT 23.18 485.64 157.32 487.35 ;
   RECT 23.18 487.35 157.32 489.06 ;
   RECT 23.18 489.06 157.32 490.77 ;
   RECT 23.18 490.77 157.32 492.48 ;
   RECT 23.18 492.48 157.32 494.19 ;
   RECT 23.18 494.19 157.32 495.9 ;
   RECT 23.18 495.9 157.32 497.61 ;
   RECT 23.18 497.61 157.32 499.32 ;
   RECT 23.18 499.32 157.32 501.03 ;
   RECT 23.18 501.03 157.32 502.74 ;
   RECT 23.18 502.74 157.32 504.45 ;
   RECT 23.18 504.45 157.32 506.16 ;
   RECT 23.18 506.16 157.32 507.87 ;
   RECT 23.18 507.87 157.32 509.58 ;
   RECT 23.18 509.58 157.32 511.29 ;
   RECT 23.18 511.29 157.32 513.0 ;
   RECT 23.18 513.0 157.32 514.71 ;
   RECT 23.18 514.71 157.32 516.42 ;
   RECT 23.18 516.42 157.32 518.13 ;
   RECT 23.18 518.13 157.32 519.84 ;
   RECT 23.18 519.84 157.32 521.55 ;
   RECT 23.18 521.55 157.32 523.26 ;
   RECT 23.18 523.26 157.32 524.97 ;
   RECT 23.18 524.97 157.32 526.68 ;
   RECT 23.18 526.68 157.32 528.39 ;
   RECT 23.18 528.39 157.32 530.1 ;
   RECT 23.18 530.1 157.32 531.81 ;
   RECT 23.18 531.81 157.32 533.52 ;
   RECT 23.18 533.52 157.32 535.23 ;
   RECT 23.18 535.23 157.32 536.94 ;
   RECT 23.18 536.94 157.32 538.65 ;
   RECT 23.18 538.65 157.32 540.36 ;
   RECT 23.18 540.36 157.32 542.07 ;
   RECT 23.18 542.07 157.32 543.78 ;
   RECT 23.18 543.78 157.32 545.49 ;
   RECT 23.18 545.49 157.32 547.2 ;
   RECT 23.18 547.2 157.32 548.91 ;
   RECT 23.18 548.91 157.32 550.62 ;
   RECT 23.18 550.62 157.32 552.33 ;
   RECT 23.18 552.33 157.32 554.04 ;
   RECT 23.18 554.04 157.32 555.75 ;
   RECT 23.18 555.75 157.32 557.46 ;
   RECT 23.18 557.46 157.32 559.17 ;
   RECT 23.18 559.17 157.32 560.88 ;
   RECT 23.18 560.88 157.32 562.59 ;
   RECT 23.18 562.59 157.32 564.3 ;
   RECT 23.18 564.3 157.32 566.01 ;
   RECT 23.18 566.01 157.32 567.72 ;
   RECT 23.18 567.72 157.32 569.43 ;
   RECT 23.18 569.43 157.32 571.14 ;
   RECT 23.18 571.14 157.32 572.85 ;
   RECT 23.18 572.85 157.32 574.56 ;
   RECT 23.18 574.56 157.32 576.27 ;
   RECT 23.18 576.27 157.32 577.98 ;
   RECT 23.18 577.98 157.32 579.69 ;
   RECT 23.18 579.69 157.32 581.4 ;
   RECT 23.18 581.4 157.32 583.11 ;
   RECT 23.18 583.11 157.32 584.82 ;
   RECT 23.18 584.82 157.32 586.53 ;
   RECT 23.18 586.53 157.32 588.24 ;
   RECT 23.18 588.24 157.32 589.95 ;
   RECT 23.18 589.95 157.32 591.66 ;
   RECT 23.18 591.66 157.32 593.37 ;
   RECT 23.18 593.37 157.32 595.08 ;
   RECT 23.18 595.08 157.32 596.79 ;
   RECT 23.18 596.79 157.32 598.5 ;
   RECT 23.18 598.5 157.32 600.21 ;
   RECT 23.18 600.21 157.32 601.92 ;
   RECT 23.18 601.92 157.32 603.63 ;
   RECT 23.18 603.63 157.32 605.34 ;
   RECT 23.18 605.34 157.32 607.05 ;
   RECT 23.18 607.05 157.32 608.76 ;
   RECT 23.18 608.76 157.32 610.47 ;
   RECT 23.18 610.47 157.32 612.18 ;
   RECT 23.18 612.18 157.32 613.89 ;
   RECT 23.18 613.89 157.32 615.6 ;
   RECT 23.18 615.6 157.32 617.31 ;
   RECT 23.18 617.31 157.32 619.02 ;
   RECT 23.18 619.02 157.32 620.73 ;
   RECT 23.18 620.73 157.32 622.44 ;
   RECT 23.18 622.44 157.32 624.15 ;
   RECT 23.18 624.15 157.32 625.86 ;
   RECT 23.18 625.86 157.32 627.57 ;
   RECT 23.18 627.57 157.32 629.28 ;
   RECT 23.18 629.28 157.32 630.99 ;
   RECT 23.18 630.99 157.32 632.7 ;
   RECT 23.18 632.7 157.32 634.41 ;
   RECT 23.18 634.41 157.32 636.12 ;
   RECT 23.18 636.12 157.32 637.83 ;
   RECT 23.18 637.83 157.32 639.54 ;
   RECT 23.18 639.54 157.32 641.25 ;
   RECT 23.18 641.25 157.32 642.96 ;
   RECT 23.18 642.96 157.32 644.67 ;
   RECT 23.18 644.67 157.32 646.38 ;
   RECT 23.18 646.38 157.32 648.09 ;
   RECT 23.18 648.09 157.32 649.8 ;
   RECT 23.18 649.8 157.32 651.51 ;
   RECT 23.18 651.51 157.32 653.22 ;
   RECT 23.18 653.22 157.32 654.93 ;
   RECT 23.18 654.93 157.32 656.64 ;
   RECT 23.18 656.64 157.32 658.35 ;
   RECT 23.18 658.35 157.32 660.06 ;
   RECT 23.18 660.06 157.32 661.77 ;
   RECT 23.18 661.77 157.32 663.48 ;
   RECT 23.18 663.48 157.32 665.19 ;
   RECT 23.18 665.19 157.32 666.9 ;
   RECT 23.18 666.9 157.32 668.61 ;
   RECT 23.18 668.61 157.32 670.32 ;
   RECT 23.18 670.32 157.32 672.03 ;
   RECT 23.18 672.03 157.32 673.74 ;
   RECT 23.18 673.74 157.32 675.45 ;
   RECT 23.18 675.45 157.32 677.16 ;
   RECT 23.18 677.16 157.32 678.87 ;
   RECT 23.18 678.87 157.32 680.58 ;
   RECT 23.18 680.58 157.32 682.29 ;
   RECT 23.18 682.29 157.32 684.0 ;
   RECT 23.18 684.0 157.32 685.71 ;
   RECT 23.18 685.71 157.32 687.42 ;
   RECT 23.18 687.42 157.32 689.13 ;
   RECT 23.18 689.13 157.32 690.84 ;
   RECT 23.18 690.84 157.32 692.55 ;
   RECT 23.18 692.55 157.32 694.26 ;
   RECT 23.18 694.26 157.32 695.97 ;
   RECT 23.18 695.97 157.32 697.68 ;
   RECT 23.18 697.68 157.32 699.39 ;
   RECT 23.18 699.39 157.32 701.1 ;
   RECT 23.18 701.1 157.32 702.81 ;
   RECT 23.18 702.81 157.32 704.52 ;
   RECT 23.18 704.52 157.32 706.23 ;
   RECT 23.18 706.23 157.32 707.94 ;
   RECT 23.18 707.94 157.32 709.65 ;
   RECT 23.18 709.65 157.32 711.36 ;
   RECT 23.18 711.36 157.32 713.07 ;
   RECT 23.18 713.07 157.32 714.78 ;
   RECT 23.18 714.78 157.32 716.49 ;
   RECT 23.18 716.49 157.32 718.2 ;
   RECT 23.18 718.2 157.32 719.91 ;
   RECT 23.18 719.91 157.32 721.62 ;
   RECT 23.18 721.62 157.32 723.33 ;
   RECT 23.18 723.33 157.32 725.04 ;
   RECT 23.18 725.04 157.32 726.75 ;
   RECT 23.18 726.75 157.32 728.46 ;
   RECT 23.18 728.46 157.32 730.17 ;
   RECT 23.18 730.17 157.32 731.88 ;
   RECT 23.18 731.88 157.32 733.59 ;
   RECT 23.18 733.59 157.32 735.3 ;
   RECT 23.18 735.3 157.32 737.01 ;
   RECT 23.18 737.01 157.32 738.72 ;
   RECT 23.18 738.72 157.32 740.43 ;
   RECT 23.18 740.43 157.32 742.14 ;
   RECT 23.18 742.14 157.32 743.85 ;
   RECT 23.18 743.85 157.32 745.56 ;
   RECT 23.18 745.56 157.32 747.27 ;
   RECT 23.18 747.27 157.32 748.98 ;
   RECT 23.18 748.98 157.32 750.69 ;
   RECT 23.18 750.69 157.32 752.4 ;
   RECT 23.18 752.4 157.32 754.11 ;
  LAYER via3 ;
   RECT 23.18 0.0 157.32 1.71 ;
   RECT 23.18 1.71 157.32 3.42 ;
   RECT 23.18 3.42 157.32 5.13 ;
   RECT 23.18 5.13 157.32 6.84 ;
   RECT 23.18 6.84 157.32 8.55 ;
   RECT 23.18 8.55 157.32 10.26 ;
   RECT 23.18 10.26 157.32 11.97 ;
   RECT 23.18 11.97 157.32 13.68 ;
   RECT 23.18 13.68 157.32 15.39 ;
   RECT 23.18 15.39 157.32 17.1 ;
   RECT 23.18 17.1 157.32 18.81 ;
   RECT 23.18 18.81 157.32 20.52 ;
   RECT 23.18 20.52 157.32 22.23 ;
   RECT 23.18 22.23 157.32 23.94 ;
   RECT 23.18 23.94 157.32 25.65 ;
   RECT 23.18 25.65 157.32 27.36 ;
   RECT 23.18 27.36 157.32 29.07 ;
   RECT 23.18 29.07 157.32 30.78 ;
   RECT 23.18 30.78 157.32 32.49 ;
   RECT 23.18 32.49 157.32 34.2 ;
   RECT 23.18 34.2 157.32 35.91 ;
   RECT 23.18 35.91 157.32 37.62 ;
   RECT 23.18 37.62 157.32 39.33 ;
   RECT 23.18 39.33 157.32 41.04 ;
   RECT 23.18 41.04 157.32 42.75 ;
   RECT 23.18 42.75 157.32 44.46 ;
   RECT 23.18 44.46 157.32 46.17 ;
   RECT 23.18 46.17 157.32 47.88 ;
   RECT 23.18 47.88 157.32 49.59 ;
   RECT 23.18 49.59 157.32 51.3 ;
   RECT 23.18 51.3 157.32 53.01 ;
   RECT 23.18 53.01 157.32 54.72 ;
   RECT 23.18 54.72 157.32 56.43 ;
   RECT 23.18 56.43 157.32 58.14 ;
   RECT 23.18 58.14 157.32 59.85 ;
   RECT 23.18 59.85 157.32 61.56 ;
   RECT 23.18 61.56 157.32 63.27 ;
   RECT 23.18 63.27 157.32 64.98 ;
   RECT 23.18 64.98 157.32 66.69 ;
   RECT 23.18 66.69 157.32 68.4 ;
   RECT 23.18 68.4 157.32 70.11 ;
   RECT 23.18 70.11 157.32 71.82 ;
   RECT 23.18 71.82 157.32 73.53 ;
   RECT 23.18 73.53 157.32 75.24 ;
   RECT 23.18 75.24 157.32 76.95 ;
   RECT 23.18 76.95 157.32 78.66 ;
   RECT 23.18 78.66 157.32 80.37 ;
   RECT 23.18 80.37 157.32 82.08 ;
   RECT 23.18 82.08 157.32 83.79 ;
   RECT 23.18 83.79 157.32 85.5 ;
   RECT 23.18 85.5 157.32 87.21 ;
   RECT 23.18 87.21 157.32 88.92 ;
   RECT 23.18 88.92 157.32 90.63 ;
   RECT 23.18 90.63 157.32 92.34 ;
   RECT 23.18 92.34 157.32 94.05 ;
   RECT 23.18 94.05 157.32 95.76 ;
   RECT 23.18 95.76 157.32 97.47 ;
   RECT 23.18 97.47 157.32 99.18 ;
   RECT 23.18 99.18 157.32 100.89 ;
   RECT 23.18 100.89 157.32 102.6 ;
   RECT 23.18 102.6 157.32 104.31 ;
   RECT 23.18 104.31 157.32 106.02 ;
   RECT 23.18 106.02 157.32 107.73 ;
   RECT 23.18 107.73 157.32 109.44 ;
   RECT 23.18 109.44 157.32 111.15 ;
   RECT 23.18 111.15 157.32 112.86 ;
   RECT 23.18 112.86 157.32 114.57 ;
   RECT 23.18 114.57 157.32 116.28 ;
   RECT 23.18 116.28 157.32 117.99 ;
   RECT 23.18 117.99 157.32 119.7 ;
   RECT 23.18 119.7 157.32 121.41 ;
   RECT 23.18 121.41 157.32 123.12 ;
   RECT 23.18 123.12 157.32 124.83 ;
   RECT 23.18 124.83 157.32 126.54 ;
   RECT 23.18 126.54 157.32 128.25 ;
   RECT 23.18 128.25 157.32 129.96 ;
   RECT 23.18 129.96 157.32 131.67 ;
   RECT 23.18 131.67 157.32 133.38 ;
   RECT 23.18 133.38 157.32 135.09 ;
   RECT 23.18 135.09 157.32 136.8 ;
   RECT 23.18 136.8 157.32 138.51 ;
   RECT 23.18 138.51 157.32 140.22 ;
   RECT 23.18 140.22 157.32 141.93 ;
   RECT 23.18 141.93 157.32 143.64 ;
   RECT 23.18 143.64 157.32 145.35 ;
   RECT 23.18 145.35 157.32 147.06 ;
   RECT 23.18 147.06 157.32 148.77 ;
   RECT 23.18 148.77 157.32 150.48 ;
   RECT 23.18 150.48 157.32 152.19 ;
   RECT 23.18 152.19 157.32 153.9 ;
   RECT 23.18 153.9 157.32 155.61 ;
   RECT 23.18 155.61 157.32 157.32 ;
   RECT 23.18 157.32 157.32 159.03 ;
   RECT 23.18 159.03 157.32 160.74 ;
   RECT 23.18 160.74 157.32 162.45 ;
   RECT 23.18 162.45 157.32 164.16 ;
   RECT 23.18 164.16 157.32 165.87 ;
   RECT 23.18 165.87 157.32 167.58 ;
   RECT 23.18 167.58 157.32 169.29 ;
   RECT 23.18 169.29 157.32 171.0 ;
   RECT 23.18 171.0 157.32 172.71 ;
   RECT 23.18 172.71 157.32 174.42 ;
   RECT 23.18 174.42 157.32 176.13 ;
   RECT 23.18 176.13 157.32 177.84 ;
   RECT 23.18 177.84 157.32 179.55 ;
   RECT 23.18 179.55 157.32 181.26 ;
   RECT 23.18 181.26 157.32 182.97 ;
   RECT 23.18 182.97 157.32 184.68 ;
   RECT 23.18 184.68 157.32 186.39 ;
   RECT 23.18 186.39 157.32 188.1 ;
   RECT 23.18 188.1 157.32 189.81 ;
   RECT 23.18 189.81 157.32 191.52 ;
   RECT 23.18 191.52 157.32 193.23 ;
   RECT 23.18 193.23 157.32 194.94 ;
   RECT 23.18 194.94 157.32 196.65 ;
   RECT 23.18 196.65 157.32 198.36 ;
   RECT 23.18 198.36 157.32 200.07 ;
   RECT 23.18 200.07 157.32 201.78 ;
   RECT 23.18 201.78 157.32 203.49 ;
   RECT 23.18 203.49 157.32 205.2 ;
   RECT 23.18 205.2 157.32 206.91 ;
   RECT 23.18 206.91 157.32 208.62 ;
   RECT 23.18 208.62 157.32 210.33 ;
   RECT 23.18 210.33 157.32 212.04 ;
   RECT 23.18 212.04 157.32 213.75 ;
   RECT 23.18 213.75 157.32 215.46 ;
   RECT 23.18 215.46 157.32 217.17 ;
   RECT 23.18 217.17 157.32 218.88 ;
   RECT 23.18 218.88 157.32 220.59 ;
   RECT 23.18 220.59 157.32 222.3 ;
   RECT 23.18 222.3 157.32 224.01 ;
   RECT 23.18 224.01 157.32 225.72 ;
   RECT 23.18 225.72 157.32 227.43 ;
   RECT 23.18 227.43 157.32 229.14 ;
   RECT 23.18 229.14 157.32 230.85 ;
   RECT 23.18 230.85 157.32 232.56 ;
   RECT 23.18 232.56 157.32 234.27 ;
   RECT 23.18 234.27 157.32 235.98 ;
   RECT 23.18 235.98 157.32 237.69 ;
   RECT 23.18 237.69 157.32 239.4 ;
   RECT 23.18 239.4 157.32 241.11 ;
   RECT 23.18 241.11 157.32 242.82 ;
   RECT 23.18 242.82 157.32 244.53 ;
   RECT 23.18 244.53 157.32 246.24 ;
   RECT 23.18 246.24 157.32 247.95 ;
   RECT 23.18 247.95 157.32 249.66 ;
   RECT 23.18 249.66 157.32 251.37 ;
   RECT 23.18 251.37 157.32 253.08 ;
   RECT 23.18 253.08 157.32 254.79 ;
   RECT 23.18 254.79 157.32 256.5 ;
   RECT 23.18 256.5 157.32 258.21 ;
   RECT 23.18 258.21 157.32 259.92 ;
   RECT 23.18 259.92 157.32 261.63 ;
   RECT 23.18 261.63 157.32 263.34 ;
   RECT 23.18 263.34 157.32 265.05 ;
   RECT 23.18 265.05 157.32 266.76 ;
   RECT 23.18 266.76 157.32 268.47 ;
   RECT 23.18 268.47 157.32 270.18 ;
   RECT 23.18 270.18 157.32 271.89 ;
   RECT 23.18 271.89 157.32 273.6 ;
   RECT 23.18 273.6 157.32 275.31 ;
   RECT 23.18 275.31 157.32 277.02 ;
   RECT 23.18 277.02 157.32 278.73 ;
   RECT 23.18 278.73 157.32 280.44 ;
   RECT 23.18 280.44 157.32 282.15 ;
   RECT 23.18 282.15 157.32 283.86 ;
   RECT 23.18 283.86 157.32 285.57 ;
   RECT 23.18 285.57 157.32 287.28 ;
   RECT 23.18 287.28 157.32 288.99 ;
   RECT 23.18 288.99 157.32 290.7 ;
   RECT 23.18 290.7 157.32 292.41 ;
   RECT 23.18 292.41 157.32 294.12 ;
   RECT 23.18 294.12 157.32 295.83 ;
   RECT 23.18 295.83 157.32 297.54 ;
   RECT 23.18 297.54 157.32 299.25 ;
   RECT 23.18 299.25 157.32 300.96 ;
   RECT 23.18 300.96 157.32 302.67 ;
   RECT 23.18 302.67 157.32 304.38 ;
   RECT 23.18 304.38 157.32 306.09 ;
   RECT 23.18 306.09 157.32 307.8 ;
   RECT 23.18 307.8 157.32 309.51 ;
   RECT 23.18 309.51 157.32 311.22 ;
   RECT 23.18 311.22 157.32 312.93 ;
   RECT 23.18 312.93 157.32 314.64 ;
   RECT 23.18 314.64 157.32 316.35 ;
   RECT 23.18 316.35 157.32 318.06 ;
   RECT 23.18 318.06 157.32 319.77 ;
   RECT 23.18 319.77 157.32 321.48 ;
   RECT 23.18 321.48 157.32 323.19 ;
   RECT 23.18 323.19 157.32 324.9 ;
   RECT 23.18 324.9 157.32 326.61 ;
   RECT 23.18 326.61 157.32 328.32 ;
   RECT 23.18 328.32 157.32 330.03 ;
   RECT 23.18 330.03 157.32 331.74 ;
   RECT 23.18 331.74 157.32 333.45 ;
   RECT 23.18 333.45 157.32 335.16 ;
   RECT 23.18 335.16 157.32 336.87 ;
   RECT 23.18 336.87 157.32 338.58 ;
   RECT 23.18 338.58 157.32 340.29 ;
   RECT 23.18 340.29 157.32 342.0 ;
   RECT 23.18 342.0 157.32 343.71 ;
   RECT 23.18 343.71 157.32 345.42 ;
   RECT 23.18 345.42 157.32 347.13 ;
   RECT 23.18 347.13 157.32 348.84 ;
   RECT 23.18 348.84 157.32 350.55 ;
   RECT 23.18 350.55 157.32 352.26 ;
   RECT 23.18 352.26 157.32 353.97 ;
   RECT 23.18 353.97 157.32 355.68 ;
   RECT 0.0 355.68 157.32 357.39 ;
   RECT 0.0 357.39 157.32 359.1 ;
   RECT 0.0 359.1 157.32 360.81 ;
   RECT 0.0 360.81 157.32 362.52 ;
   RECT 0.0 362.52 157.32 364.23 ;
   RECT 0.0 364.23 157.32 365.94 ;
   RECT 0.0 365.94 157.32 367.65 ;
   RECT 0.0 367.65 157.32 369.36 ;
   RECT 0.0 369.36 157.32 371.07 ;
   RECT 0.0 371.07 157.32 372.78 ;
   RECT 0.0 372.78 157.32 374.49 ;
   RECT 0.0 374.49 157.32 376.2 ;
   RECT 0.0 376.2 157.32 377.91 ;
   RECT 0.0 377.91 157.32 379.62 ;
   RECT 0.0 379.62 157.32 381.33 ;
   RECT 0.0 381.33 157.32 383.04 ;
   RECT 0.0 383.04 157.32 384.75 ;
   RECT 23.18 384.75 157.32 386.46 ;
   RECT 23.18 386.46 157.32 388.17 ;
   RECT 23.18 388.17 157.32 389.88 ;
   RECT 23.18 389.88 157.32 391.59 ;
   RECT 23.18 391.59 157.32 393.3 ;
   RECT 23.18 393.3 157.32 395.01 ;
   RECT 23.18 395.01 157.32 396.72 ;
   RECT 23.18 396.72 157.32 398.43 ;
   RECT 23.18 398.43 157.32 400.14 ;
   RECT 23.18 400.14 157.32 401.85 ;
   RECT 23.18 401.85 157.32 403.56 ;
   RECT 23.18 403.56 157.32 405.27 ;
   RECT 23.18 405.27 157.32 406.98 ;
   RECT 23.18 406.98 157.32 408.69 ;
   RECT 23.18 408.69 157.32 410.4 ;
   RECT 23.18 410.4 157.32 412.11 ;
   RECT 23.18 412.11 157.32 413.82 ;
   RECT 23.18 413.82 157.32 415.53 ;
   RECT 23.18 415.53 157.32 417.24 ;
   RECT 23.18 417.24 157.32 418.95 ;
   RECT 23.18 418.95 157.32 420.66 ;
   RECT 23.18 420.66 157.32 422.37 ;
   RECT 23.18 422.37 157.32 424.08 ;
   RECT 23.18 424.08 157.32 425.79 ;
   RECT 23.18 425.79 157.32 427.5 ;
   RECT 23.18 427.5 157.32 429.21 ;
   RECT 23.18 429.21 157.32 430.92 ;
   RECT 23.18 430.92 157.32 432.63 ;
   RECT 23.18 432.63 157.32 434.34 ;
   RECT 23.18 434.34 157.32 436.05 ;
   RECT 23.18 436.05 157.32 437.76 ;
   RECT 23.18 437.76 157.32 439.47 ;
   RECT 23.18 439.47 157.32 441.18 ;
   RECT 23.18 441.18 157.32 442.89 ;
   RECT 23.18 442.89 157.32 444.6 ;
   RECT 23.18 444.6 157.32 446.31 ;
   RECT 23.18 446.31 157.32 448.02 ;
   RECT 23.18 448.02 157.32 449.73 ;
   RECT 23.18 449.73 157.32 451.44 ;
   RECT 23.18 451.44 157.32 453.15 ;
   RECT 23.18 453.15 157.32 454.86 ;
   RECT 23.18 454.86 157.32 456.57 ;
   RECT 23.18 456.57 157.32 458.28 ;
   RECT 23.18 458.28 157.32 459.99 ;
   RECT 23.18 459.99 157.32 461.7 ;
   RECT 23.18 461.7 157.32 463.41 ;
   RECT 23.18 463.41 157.32 465.12 ;
   RECT 23.18 465.12 157.32 466.83 ;
   RECT 23.18 466.83 157.32 468.54 ;
   RECT 23.18 468.54 157.32 470.25 ;
   RECT 23.18 470.25 157.32 471.96 ;
   RECT 23.18 471.96 157.32 473.67 ;
   RECT 23.18 473.67 157.32 475.38 ;
   RECT 23.18 475.38 157.32 477.09 ;
   RECT 23.18 477.09 157.32 478.8 ;
   RECT 23.18 478.8 157.32 480.51 ;
   RECT 23.18 480.51 157.32 482.22 ;
   RECT 23.18 482.22 157.32 483.93 ;
   RECT 23.18 483.93 157.32 485.64 ;
   RECT 23.18 485.64 157.32 487.35 ;
   RECT 23.18 487.35 157.32 489.06 ;
   RECT 23.18 489.06 157.32 490.77 ;
   RECT 23.18 490.77 157.32 492.48 ;
   RECT 23.18 492.48 157.32 494.19 ;
   RECT 23.18 494.19 157.32 495.9 ;
   RECT 23.18 495.9 157.32 497.61 ;
   RECT 23.18 497.61 157.32 499.32 ;
   RECT 23.18 499.32 157.32 501.03 ;
   RECT 23.18 501.03 157.32 502.74 ;
   RECT 23.18 502.74 157.32 504.45 ;
   RECT 23.18 504.45 157.32 506.16 ;
   RECT 23.18 506.16 157.32 507.87 ;
   RECT 23.18 507.87 157.32 509.58 ;
   RECT 23.18 509.58 157.32 511.29 ;
   RECT 23.18 511.29 157.32 513.0 ;
   RECT 23.18 513.0 157.32 514.71 ;
   RECT 23.18 514.71 157.32 516.42 ;
   RECT 23.18 516.42 157.32 518.13 ;
   RECT 23.18 518.13 157.32 519.84 ;
   RECT 23.18 519.84 157.32 521.55 ;
   RECT 23.18 521.55 157.32 523.26 ;
   RECT 23.18 523.26 157.32 524.97 ;
   RECT 23.18 524.97 157.32 526.68 ;
   RECT 23.18 526.68 157.32 528.39 ;
   RECT 23.18 528.39 157.32 530.1 ;
   RECT 23.18 530.1 157.32 531.81 ;
   RECT 23.18 531.81 157.32 533.52 ;
   RECT 23.18 533.52 157.32 535.23 ;
   RECT 23.18 535.23 157.32 536.94 ;
   RECT 23.18 536.94 157.32 538.65 ;
   RECT 23.18 538.65 157.32 540.36 ;
   RECT 23.18 540.36 157.32 542.07 ;
   RECT 23.18 542.07 157.32 543.78 ;
   RECT 23.18 543.78 157.32 545.49 ;
   RECT 23.18 545.49 157.32 547.2 ;
   RECT 23.18 547.2 157.32 548.91 ;
   RECT 23.18 548.91 157.32 550.62 ;
   RECT 23.18 550.62 157.32 552.33 ;
   RECT 23.18 552.33 157.32 554.04 ;
   RECT 23.18 554.04 157.32 555.75 ;
   RECT 23.18 555.75 157.32 557.46 ;
   RECT 23.18 557.46 157.32 559.17 ;
   RECT 23.18 559.17 157.32 560.88 ;
   RECT 23.18 560.88 157.32 562.59 ;
   RECT 23.18 562.59 157.32 564.3 ;
   RECT 23.18 564.3 157.32 566.01 ;
   RECT 23.18 566.01 157.32 567.72 ;
   RECT 23.18 567.72 157.32 569.43 ;
   RECT 23.18 569.43 157.32 571.14 ;
   RECT 23.18 571.14 157.32 572.85 ;
   RECT 23.18 572.85 157.32 574.56 ;
   RECT 23.18 574.56 157.32 576.27 ;
   RECT 23.18 576.27 157.32 577.98 ;
   RECT 23.18 577.98 157.32 579.69 ;
   RECT 23.18 579.69 157.32 581.4 ;
   RECT 23.18 581.4 157.32 583.11 ;
   RECT 23.18 583.11 157.32 584.82 ;
   RECT 23.18 584.82 157.32 586.53 ;
   RECT 23.18 586.53 157.32 588.24 ;
   RECT 23.18 588.24 157.32 589.95 ;
   RECT 23.18 589.95 157.32 591.66 ;
   RECT 23.18 591.66 157.32 593.37 ;
   RECT 23.18 593.37 157.32 595.08 ;
   RECT 23.18 595.08 157.32 596.79 ;
   RECT 23.18 596.79 157.32 598.5 ;
   RECT 23.18 598.5 157.32 600.21 ;
   RECT 23.18 600.21 157.32 601.92 ;
   RECT 23.18 601.92 157.32 603.63 ;
   RECT 23.18 603.63 157.32 605.34 ;
   RECT 23.18 605.34 157.32 607.05 ;
   RECT 23.18 607.05 157.32 608.76 ;
   RECT 23.18 608.76 157.32 610.47 ;
   RECT 23.18 610.47 157.32 612.18 ;
   RECT 23.18 612.18 157.32 613.89 ;
   RECT 23.18 613.89 157.32 615.6 ;
   RECT 23.18 615.6 157.32 617.31 ;
   RECT 23.18 617.31 157.32 619.02 ;
   RECT 23.18 619.02 157.32 620.73 ;
   RECT 23.18 620.73 157.32 622.44 ;
   RECT 23.18 622.44 157.32 624.15 ;
   RECT 23.18 624.15 157.32 625.86 ;
   RECT 23.18 625.86 157.32 627.57 ;
   RECT 23.18 627.57 157.32 629.28 ;
   RECT 23.18 629.28 157.32 630.99 ;
   RECT 23.18 630.99 157.32 632.7 ;
   RECT 23.18 632.7 157.32 634.41 ;
   RECT 23.18 634.41 157.32 636.12 ;
   RECT 23.18 636.12 157.32 637.83 ;
   RECT 23.18 637.83 157.32 639.54 ;
   RECT 23.18 639.54 157.32 641.25 ;
   RECT 23.18 641.25 157.32 642.96 ;
   RECT 23.18 642.96 157.32 644.67 ;
   RECT 23.18 644.67 157.32 646.38 ;
   RECT 23.18 646.38 157.32 648.09 ;
   RECT 23.18 648.09 157.32 649.8 ;
   RECT 23.18 649.8 157.32 651.51 ;
   RECT 23.18 651.51 157.32 653.22 ;
   RECT 23.18 653.22 157.32 654.93 ;
   RECT 23.18 654.93 157.32 656.64 ;
   RECT 23.18 656.64 157.32 658.35 ;
   RECT 23.18 658.35 157.32 660.06 ;
   RECT 23.18 660.06 157.32 661.77 ;
   RECT 23.18 661.77 157.32 663.48 ;
   RECT 23.18 663.48 157.32 665.19 ;
   RECT 23.18 665.19 157.32 666.9 ;
   RECT 23.18 666.9 157.32 668.61 ;
   RECT 23.18 668.61 157.32 670.32 ;
   RECT 23.18 670.32 157.32 672.03 ;
   RECT 23.18 672.03 157.32 673.74 ;
   RECT 23.18 673.74 157.32 675.45 ;
   RECT 23.18 675.45 157.32 677.16 ;
   RECT 23.18 677.16 157.32 678.87 ;
   RECT 23.18 678.87 157.32 680.58 ;
   RECT 23.18 680.58 157.32 682.29 ;
   RECT 23.18 682.29 157.32 684.0 ;
   RECT 23.18 684.0 157.32 685.71 ;
   RECT 23.18 685.71 157.32 687.42 ;
   RECT 23.18 687.42 157.32 689.13 ;
   RECT 23.18 689.13 157.32 690.84 ;
   RECT 23.18 690.84 157.32 692.55 ;
   RECT 23.18 692.55 157.32 694.26 ;
   RECT 23.18 694.26 157.32 695.97 ;
   RECT 23.18 695.97 157.32 697.68 ;
   RECT 23.18 697.68 157.32 699.39 ;
   RECT 23.18 699.39 157.32 701.1 ;
   RECT 23.18 701.1 157.32 702.81 ;
   RECT 23.18 702.81 157.32 704.52 ;
   RECT 23.18 704.52 157.32 706.23 ;
   RECT 23.18 706.23 157.32 707.94 ;
   RECT 23.18 707.94 157.32 709.65 ;
   RECT 23.18 709.65 157.32 711.36 ;
   RECT 23.18 711.36 157.32 713.07 ;
   RECT 23.18 713.07 157.32 714.78 ;
   RECT 23.18 714.78 157.32 716.49 ;
   RECT 23.18 716.49 157.32 718.2 ;
   RECT 23.18 718.2 157.32 719.91 ;
   RECT 23.18 719.91 157.32 721.62 ;
   RECT 23.18 721.62 157.32 723.33 ;
   RECT 23.18 723.33 157.32 725.04 ;
   RECT 23.18 725.04 157.32 726.75 ;
   RECT 23.18 726.75 157.32 728.46 ;
   RECT 23.18 728.46 157.32 730.17 ;
   RECT 23.18 730.17 157.32 731.88 ;
   RECT 23.18 731.88 157.32 733.59 ;
   RECT 23.18 733.59 157.32 735.3 ;
   RECT 23.18 735.3 157.32 737.01 ;
   RECT 23.18 737.01 157.32 738.72 ;
   RECT 23.18 738.72 157.32 740.43 ;
   RECT 23.18 740.43 157.32 742.14 ;
   RECT 23.18 742.14 157.32 743.85 ;
   RECT 23.18 743.85 157.32 745.56 ;
   RECT 23.18 745.56 157.32 747.27 ;
   RECT 23.18 747.27 157.32 748.98 ;
   RECT 23.18 748.98 157.32 750.69 ;
   RECT 23.18 750.69 157.32 752.4 ;
   RECT 23.18 752.4 157.32 754.11 ;
  LAYER metal4 ;
   RECT 23.18 0.0 157.32 1.71 ;
   RECT 23.18 1.71 157.32 3.42 ;
   RECT 23.18 3.42 157.32 5.13 ;
   RECT 23.18 5.13 157.32 6.84 ;
   RECT 23.18 6.84 157.32 8.55 ;
   RECT 23.18 8.55 157.32 10.26 ;
   RECT 23.18 10.26 157.32 11.97 ;
   RECT 23.18 11.97 157.32 13.68 ;
   RECT 23.18 13.68 157.32 15.39 ;
   RECT 23.18 15.39 157.32 17.1 ;
   RECT 23.18 17.1 157.32 18.81 ;
   RECT 23.18 18.81 157.32 20.52 ;
   RECT 23.18 20.52 157.32 22.23 ;
   RECT 23.18 22.23 157.32 23.94 ;
   RECT 23.18 23.94 157.32 25.65 ;
   RECT 23.18 25.65 157.32 27.36 ;
   RECT 23.18 27.36 157.32 29.07 ;
   RECT 23.18 29.07 157.32 30.78 ;
   RECT 23.18 30.78 157.32 32.49 ;
   RECT 23.18 32.49 157.32 34.2 ;
   RECT 23.18 34.2 157.32 35.91 ;
   RECT 23.18 35.91 157.32 37.62 ;
   RECT 23.18 37.62 157.32 39.33 ;
   RECT 23.18 39.33 157.32 41.04 ;
   RECT 23.18 41.04 157.32 42.75 ;
   RECT 23.18 42.75 157.32 44.46 ;
   RECT 23.18 44.46 157.32 46.17 ;
   RECT 23.18 46.17 157.32 47.88 ;
   RECT 23.18 47.88 157.32 49.59 ;
   RECT 23.18 49.59 157.32 51.3 ;
   RECT 23.18 51.3 157.32 53.01 ;
   RECT 23.18 53.01 157.32 54.72 ;
   RECT 23.18 54.72 157.32 56.43 ;
   RECT 23.18 56.43 157.32 58.14 ;
   RECT 23.18 58.14 157.32 59.85 ;
   RECT 23.18 59.85 157.32 61.56 ;
   RECT 23.18 61.56 157.32 63.27 ;
   RECT 23.18 63.27 157.32 64.98 ;
   RECT 23.18 64.98 157.32 66.69 ;
   RECT 23.18 66.69 157.32 68.4 ;
   RECT 23.18 68.4 157.32 70.11 ;
   RECT 23.18 70.11 157.32 71.82 ;
   RECT 23.18 71.82 157.32 73.53 ;
   RECT 23.18 73.53 157.32 75.24 ;
   RECT 23.18 75.24 157.32 76.95 ;
   RECT 23.18 76.95 157.32 78.66 ;
   RECT 23.18 78.66 157.32 80.37 ;
   RECT 23.18 80.37 157.32 82.08 ;
   RECT 23.18 82.08 157.32 83.79 ;
   RECT 23.18 83.79 157.32 85.5 ;
   RECT 23.18 85.5 157.32 87.21 ;
   RECT 23.18 87.21 157.32 88.92 ;
   RECT 23.18 88.92 157.32 90.63 ;
   RECT 23.18 90.63 157.32 92.34 ;
   RECT 23.18 92.34 157.32 94.05 ;
   RECT 23.18 94.05 157.32 95.76 ;
   RECT 23.18 95.76 157.32 97.47 ;
   RECT 23.18 97.47 157.32 99.18 ;
   RECT 23.18 99.18 157.32 100.89 ;
   RECT 23.18 100.89 157.32 102.6 ;
   RECT 23.18 102.6 157.32 104.31 ;
   RECT 23.18 104.31 157.32 106.02 ;
   RECT 23.18 106.02 157.32 107.73 ;
   RECT 23.18 107.73 157.32 109.44 ;
   RECT 23.18 109.44 157.32 111.15 ;
   RECT 23.18 111.15 157.32 112.86 ;
   RECT 23.18 112.86 157.32 114.57 ;
   RECT 23.18 114.57 157.32 116.28 ;
   RECT 23.18 116.28 157.32 117.99 ;
   RECT 23.18 117.99 157.32 119.7 ;
   RECT 23.18 119.7 157.32 121.41 ;
   RECT 23.18 121.41 157.32 123.12 ;
   RECT 23.18 123.12 157.32 124.83 ;
   RECT 23.18 124.83 157.32 126.54 ;
   RECT 23.18 126.54 157.32 128.25 ;
   RECT 23.18 128.25 157.32 129.96 ;
   RECT 23.18 129.96 157.32 131.67 ;
   RECT 23.18 131.67 157.32 133.38 ;
   RECT 23.18 133.38 157.32 135.09 ;
   RECT 23.18 135.09 157.32 136.8 ;
   RECT 23.18 136.8 157.32 138.51 ;
   RECT 23.18 138.51 157.32 140.22 ;
   RECT 23.18 140.22 157.32 141.93 ;
   RECT 23.18 141.93 157.32 143.64 ;
   RECT 23.18 143.64 157.32 145.35 ;
   RECT 23.18 145.35 157.32 147.06 ;
   RECT 23.18 147.06 157.32 148.77 ;
   RECT 23.18 148.77 157.32 150.48 ;
   RECT 23.18 150.48 157.32 152.19 ;
   RECT 23.18 152.19 157.32 153.9 ;
   RECT 23.18 153.9 157.32 155.61 ;
   RECT 23.18 155.61 157.32 157.32 ;
   RECT 23.18 157.32 157.32 159.03 ;
   RECT 23.18 159.03 157.32 160.74 ;
   RECT 23.18 160.74 157.32 162.45 ;
   RECT 23.18 162.45 157.32 164.16 ;
   RECT 23.18 164.16 157.32 165.87 ;
   RECT 23.18 165.87 157.32 167.58 ;
   RECT 23.18 167.58 157.32 169.29 ;
   RECT 23.18 169.29 157.32 171.0 ;
   RECT 23.18 171.0 157.32 172.71 ;
   RECT 23.18 172.71 157.32 174.42 ;
   RECT 23.18 174.42 157.32 176.13 ;
   RECT 23.18 176.13 157.32 177.84 ;
   RECT 23.18 177.84 157.32 179.55 ;
   RECT 23.18 179.55 157.32 181.26 ;
   RECT 23.18 181.26 157.32 182.97 ;
   RECT 23.18 182.97 157.32 184.68 ;
   RECT 23.18 184.68 157.32 186.39 ;
   RECT 23.18 186.39 157.32 188.1 ;
   RECT 23.18 188.1 157.32 189.81 ;
   RECT 23.18 189.81 157.32 191.52 ;
   RECT 23.18 191.52 157.32 193.23 ;
   RECT 23.18 193.23 157.32 194.94 ;
   RECT 23.18 194.94 157.32 196.65 ;
   RECT 23.18 196.65 157.32 198.36 ;
   RECT 23.18 198.36 157.32 200.07 ;
   RECT 23.18 200.07 157.32 201.78 ;
   RECT 23.18 201.78 157.32 203.49 ;
   RECT 23.18 203.49 157.32 205.2 ;
   RECT 23.18 205.2 157.32 206.91 ;
   RECT 23.18 206.91 157.32 208.62 ;
   RECT 23.18 208.62 157.32 210.33 ;
   RECT 23.18 210.33 157.32 212.04 ;
   RECT 23.18 212.04 157.32 213.75 ;
   RECT 23.18 213.75 157.32 215.46 ;
   RECT 23.18 215.46 157.32 217.17 ;
   RECT 23.18 217.17 157.32 218.88 ;
   RECT 23.18 218.88 157.32 220.59 ;
   RECT 23.18 220.59 157.32 222.3 ;
   RECT 23.18 222.3 157.32 224.01 ;
   RECT 23.18 224.01 157.32 225.72 ;
   RECT 23.18 225.72 157.32 227.43 ;
   RECT 23.18 227.43 157.32 229.14 ;
   RECT 23.18 229.14 157.32 230.85 ;
   RECT 23.18 230.85 157.32 232.56 ;
   RECT 23.18 232.56 157.32 234.27 ;
   RECT 23.18 234.27 157.32 235.98 ;
   RECT 23.18 235.98 157.32 237.69 ;
   RECT 23.18 237.69 157.32 239.4 ;
   RECT 23.18 239.4 157.32 241.11 ;
   RECT 23.18 241.11 157.32 242.82 ;
   RECT 23.18 242.82 157.32 244.53 ;
   RECT 23.18 244.53 157.32 246.24 ;
   RECT 23.18 246.24 157.32 247.95 ;
   RECT 23.18 247.95 157.32 249.66 ;
   RECT 23.18 249.66 157.32 251.37 ;
   RECT 23.18 251.37 157.32 253.08 ;
   RECT 23.18 253.08 157.32 254.79 ;
   RECT 23.18 254.79 157.32 256.5 ;
   RECT 23.18 256.5 157.32 258.21 ;
   RECT 23.18 258.21 157.32 259.92 ;
   RECT 23.18 259.92 157.32 261.63 ;
   RECT 23.18 261.63 157.32 263.34 ;
   RECT 23.18 263.34 157.32 265.05 ;
   RECT 23.18 265.05 157.32 266.76 ;
   RECT 23.18 266.76 157.32 268.47 ;
   RECT 23.18 268.47 157.32 270.18 ;
   RECT 23.18 270.18 157.32 271.89 ;
   RECT 23.18 271.89 157.32 273.6 ;
   RECT 23.18 273.6 157.32 275.31 ;
   RECT 23.18 275.31 157.32 277.02 ;
   RECT 23.18 277.02 157.32 278.73 ;
   RECT 23.18 278.73 157.32 280.44 ;
   RECT 23.18 280.44 157.32 282.15 ;
   RECT 23.18 282.15 157.32 283.86 ;
   RECT 23.18 283.86 157.32 285.57 ;
   RECT 23.18 285.57 157.32 287.28 ;
   RECT 23.18 287.28 157.32 288.99 ;
   RECT 23.18 288.99 157.32 290.7 ;
   RECT 23.18 290.7 157.32 292.41 ;
   RECT 23.18 292.41 157.32 294.12 ;
   RECT 23.18 294.12 157.32 295.83 ;
   RECT 23.18 295.83 157.32 297.54 ;
   RECT 23.18 297.54 157.32 299.25 ;
   RECT 23.18 299.25 157.32 300.96 ;
   RECT 23.18 300.96 157.32 302.67 ;
   RECT 23.18 302.67 157.32 304.38 ;
   RECT 23.18 304.38 157.32 306.09 ;
   RECT 23.18 306.09 157.32 307.8 ;
   RECT 23.18 307.8 157.32 309.51 ;
   RECT 23.18 309.51 157.32 311.22 ;
   RECT 23.18 311.22 157.32 312.93 ;
   RECT 23.18 312.93 157.32 314.64 ;
   RECT 23.18 314.64 157.32 316.35 ;
   RECT 23.18 316.35 157.32 318.06 ;
   RECT 23.18 318.06 157.32 319.77 ;
   RECT 23.18 319.77 157.32 321.48 ;
   RECT 23.18 321.48 157.32 323.19 ;
   RECT 23.18 323.19 157.32 324.9 ;
   RECT 23.18 324.9 157.32 326.61 ;
   RECT 23.18 326.61 157.32 328.32 ;
   RECT 23.18 328.32 157.32 330.03 ;
   RECT 23.18 330.03 157.32 331.74 ;
   RECT 23.18 331.74 157.32 333.45 ;
   RECT 23.18 333.45 157.32 335.16 ;
   RECT 23.18 335.16 157.32 336.87 ;
   RECT 23.18 336.87 157.32 338.58 ;
   RECT 23.18 338.58 157.32 340.29 ;
   RECT 23.18 340.29 157.32 342.0 ;
   RECT 23.18 342.0 157.32 343.71 ;
   RECT 23.18 343.71 157.32 345.42 ;
   RECT 23.18 345.42 157.32 347.13 ;
   RECT 23.18 347.13 157.32 348.84 ;
   RECT 23.18 348.84 157.32 350.55 ;
   RECT 23.18 350.55 157.32 352.26 ;
   RECT 23.18 352.26 157.32 353.97 ;
   RECT 23.18 353.97 157.32 355.68 ;
   RECT 0.0 355.68 157.32 357.39 ;
   RECT 0.0 357.39 157.32 359.1 ;
   RECT 0.0 359.1 157.32 360.81 ;
   RECT 0.0 360.81 157.32 362.52 ;
   RECT 0.0 362.52 157.32 364.23 ;
   RECT 0.0 364.23 157.32 365.94 ;
   RECT 0.0 365.94 157.32 367.65 ;
   RECT 0.0 367.65 157.32 369.36 ;
   RECT 0.0 369.36 157.32 371.07 ;
   RECT 0.0 371.07 157.32 372.78 ;
   RECT 0.0 372.78 157.32 374.49 ;
   RECT 0.0 374.49 157.32 376.2 ;
   RECT 0.0 376.2 157.32 377.91 ;
   RECT 0.0 377.91 157.32 379.62 ;
   RECT 0.0 379.62 157.32 381.33 ;
   RECT 0.0 381.33 157.32 383.04 ;
   RECT 0.0 383.04 157.32 384.75 ;
   RECT 23.18 384.75 157.32 386.46 ;
   RECT 23.18 386.46 157.32 388.17 ;
   RECT 23.18 388.17 157.32 389.88 ;
   RECT 23.18 389.88 157.32 391.59 ;
   RECT 23.18 391.59 157.32 393.3 ;
   RECT 23.18 393.3 157.32 395.01 ;
   RECT 23.18 395.01 157.32 396.72 ;
   RECT 23.18 396.72 157.32 398.43 ;
   RECT 23.18 398.43 157.32 400.14 ;
   RECT 23.18 400.14 157.32 401.85 ;
   RECT 23.18 401.85 157.32 403.56 ;
   RECT 23.18 403.56 157.32 405.27 ;
   RECT 23.18 405.27 157.32 406.98 ;
   RECT 23.18 406.98 157.32 408.69 ;
   RECT 23.18 408.69 157.32 410.4 ;
   RECT 23.18 410.4 157.32 412.11 ;
   RECT 23.18 412.11 157.32 413.82 ;
   RECT 23.18 413.82 157.32 415.53 ;
   RECT 23.18 415.53 157.32 417.24 ;
   RECT 23.18 417.24 157.32 418.95 ;
   RECT 23.18 418.95 157.32 420.66 ;
   RECT 23.18 420.66 157.32 422.37 ;
   RECT 23.18 422.37 157.32 424.08 ;
   RECT 23.18 424.08 157.32 425.79 ;
   RECT 23.18 425.79 157.32 427.5 ;
   RECT 23.18 427.5 157.32 429.21 ;
   RECT 23.18 429.21 157.32 430.92 ;
   RECT 23.18 430.92 157.32 432.63 ;
   RECT 23.18 432.63 157.32 434.34 ;
   RECT 23.18 434.34 157.32 436.05 ;
   RECT 23.18 436.05 157.32 437.76 ;
   RECT 23.18 437.76 157.32 439.47 ;
   RECT 23.18 439.47 157.32 441.18 ;
   RECT 23.18 441.18 157.32 442.89 ;
   RECT 23.18 442.89 157.32 444.6 ;
   RECT 23.18 444.6 157.32 446.31 ;
   RECT 23.18 446.31 157.32 448.02 ;
   RECT 23.18 448.02 157.32 449.73 ;
   RECT 23.18 449.73 157.32 451.44 ;
   RECT 23.18 451.44 157.32 453.15 ;
   RECT 23.18 453.15 157.32 454.86 ;
   RECT 23.18 454.86 157.32 456.57 ;
   RECT 23.18 456.57 157.32 458.28 ;
   RECT 23.18 458.28 157.32 459.99 ;
   RECT 23.18 459.99 157.32 461.7 ;
   RECT 23.18 461.7 157.32 463.41 ;
   RECT 23.18 463.41 157.32 465.12 ;
   RECT 23.18 465.12 157.32 466.83 ;
   RECT 23.18 466.83 157.32 468.54 ;
   RECT 23.18 468.54 157.32 470.25 ;
   RECT 23.18 470.25 157.32 471.96 ;
   RECT 23.18 471.96 157.32 473.67 ;
   RECT 23.18 473.67 157.32 475.38 ;
   RECT 23.18 475.38 157.32 477.09 ;
   RECT 23.18 477.09 157.32 478.8 ;
   RECT 23.18 478.8 157.32 480.51 ;
   RECT 23.18 480.51 157.32 482.22 ;
   RECT 23.18 482.22 157.32 483.93 ;
   RECT 23.18 483.93 157.32 485.64 ;
   RECT 23.18 485.64 157.32 487.35 ;
   RECT 23.18 487.35 157.32 489.06 ;
   RECT 23.18 489.06 157.32 490.77 ;
   RECT 23.18 490.77 157.32 492.48 ;
   RECT 23.18 492.48 157.32 494.19 ;
   RECT 23.18 494.19 157.32 495.9 ;
   RECT 23.18 495.9 157.32 497.61 ;
   RECT 23.18 497.61 157.32 499.32 ;
   RECT 23.18 499.32 157.32 501.03 ;
   RECT 23.18 501.03 157.32 502.74 ;
   RECT 23.18 502.74 157.32 504.45 ;
   RECT 23.18 504.45 157.32 506.16 ;
   RECT 23.18 506.16 157.32 507.87 ;
   RECT 23.18 507.87 157.32 509.58 ;
   RECT 23.18 509.58 157.32 511.29 ;
   RECT 23.18 511.29 157.32 513.0 ;
   RECT 23.18 513.0 157.32 514.71 ;
   RECT 23.18 514.71 157.32 516.42 ;
   RECT 23.18 516.42 157.32 518.13 ;
   RECT 23.18 518.13 157.32 519.84 ;
   RECT 23.18 519.84 157.32 521.55 ;
   RECT 23.18 521.55 157.32 523.26 ;
   RECT 23.18 523.26 157.32 524.97 ;
   RECT 23.18 524.97 157.32 526.68 ;
   RECT 23.18 526.68 157.32 528.39 ;
   RECT 23.18 528.39 157.32 530.1 ;
   RECT 23.18 530.1 157.32 531.81 ;
   RECT 23.18 531.81 157.32 533.52 ;
   RECT 23.18 533.52 157.32 535.23 ;
   RECT 23.18 535.23 157.32 536.94 ;
   RECT 23.18 536.94 157.32 538.65 ;
   RECT 23.18 538.65 157.32 540.36 ;
   RECT 23.18 540.36 157.32 542.07 ;
   RECT 23.18 542.07 157.32 543.78 ;
   RECT 23.18 543.78 157.32 545.49 ;
   RECT 23.18 545.49 157.32 547.2 ;
   RECT 23.18 547.2 157.32 548.91 ;
   RECT 23.18 548.91 157.32 550.62 ;
   RECT 23.18 550.62 157.32 552.33 ;
   RECT 23.18 552.33 157.32 554.04 ;
   RECT 23.18 554.04 157.32 555.75 ;
   RECT 23.18 555.75 157.32 557.46 ;
   RECT 23.18 557.46 157.32 559.17 ;
   RECT 23.18 559.17 157.32 560.88 ;
   RECT 23.18 560.88 157.32 562.59 ;
   RECT 23.18 562.59 157.32 564.3 ;
   RECT 23.18 564.3 157.32 566.01 ;
   RECT 23.18 566.01 157.32 567.72 ;
   RECT 23.18 567.72 157.32 569.43 ;
   RECT 23.18 569.43 157.32 571.14 ;
   RECT 23.18 571.14 157.32 572.85 ;
   RECT 23.18 572.85 157.32 574.56 ;
   RECT 23.18 574.56 157.32 576.27 ;
   RECT 23.18 576.27 157.32 577.98 ;
   RECT 23.18 577.98 157.32 579.69 ;
   RECT 23.18 579.69 157.32 581.4 ;
   RECT 23.18 581.4 157.32 583.11 ;
   RECT 23.18 583.11 157.32 584.82 ;
   RECT 23.18 584.82 157.32 586.53 ;
   RECT 23.18 586.53 157.32 588.24 ;
   RECT 23.18 588.24 157.32 589.95 ;
   RECT 23.18 589.95 157.32 591.66 ;
   RECT 23.18 591.66 157.32 593.37 ;
   RECT 23.18 593.37 157.32 595.08 ;
   RECT 23.18 595.08 157.32 596.79 ;
   RECT 23.18 596.79 157.32 598.5 ;
   RECT 23.18 598.5 157.32 600.21 ;
   RECT 23.18 600.21 157.32 601.92 ;
   RECT 23.18 601.92 157.32 603.63 ;
   RECT 23.18 603.63 157.32 605.34 ;
   RECT 23.18 605.34 157.32 607.05 ;
   RECT 23.18 607.05 157.32 608.76 ;
   RECT 23.18 608.76 157.32 610.47 ;
   RECT 23.18 610.47 157.32 612.18 ;
   RECT 23.18 612.18 157.32 613.89 ;
   RECT 23.18 613.89 157.32 615.6 ;
   RECT 23.18 615.6 157.32 617.31 ;
   RECT 23.18 617.31 157.32 619.02 ;
   RECT 23.18 619.02 157.32 620.73 ;
   RECT 23.18 620.73 157.32 622.44 ;
   RECT 23.18 622.44 157.32 624.15 ;
   RECT 23.18 624.15 157.32 625.86 ;
   RECT 23.18 625.86 157.32 627.57 ;
   RECT 23.18 627.57 157.32 629.28 ;
   RECT 23.18 629.28 157.32 630.99 ;
   RECT 23.18 630.99 157.32 632.7 ;
   RECT 23.18 632.7 157.32 634.41 ;
   RECT 23.18 634.41 157.32 636.12 ;
   RECT 23.18 636.12 157.32 637.83 ;
   RECT 23.18 637.83 157.32 639.54 ;
   RECT 23.18 639.54 157.32 641.25 ;
   RECT 23.18 641.25 157.32 642.96 ;
   RECT 23.18 642.96 157.32 644.67 ;
   RECT 23.18 644.67 157.32 646.38 ;
   RECT 23.18 646.38 157.32 648.09 ;
   RECT 23.18 648.09 157.32 649.8 ;
   RECT 23.18 649.8 157.32 651.51 ;
   RECT 23.18 651.51 157.32 653.22 ;
   RECT 23.18 653.22 157.32 654.93 ;
   RECT 23.18 654.93 157.32 656.64 ;
   RECT 23.18 656.64 157.32 658.35 ;
   RECT 23.18 658.35 157.32 660.06 ;
   RECT 23.18 660.06 157.32 661.77 ;
   RECT 23.18 661.77 157.32 663.48 ;
   RECT 23.18 663.48 157.32 665.19 ;
   RECT 23.18 665.19 157.32 666.9 ;
   RECT 23.18 666.9 157.32 668.61 ;
   RECT 23.18 668.61 157.32 670.32 ;
   RECT 23.18 670.32 157.32 672.03 ;
   RECT 23.18 672.03 157.32 673.74 ;
   RECT 23.18 673.74 157.32 675.45 ;
   RECT 23.18 675.45 157.32 677.16 ;
   RECT 23.18 677.16 157.32 678.87 ;
   RECT 23.18 678.87 157.32 680.58 ;
   RECT 23.18 680.58 157.32 682.29 ;
   RECT 23.18 682.29 157.32 684.0 ;
   RECT 23.18 684.0 157.32 685.71 ;
   RECT 23.18 685.71 157.32 687.42 ;
   RECT 23.18 687.42 157.32 689.13 ;
   RECT 23.18 689.13 157.32 690.84 ;
   RECT 23.18 690.84 157.32 692.55 ;
   RECT 23.18 692.55 157.32 694.26 ;
   RECT 23.18 694.26 157.32 695.97 ;
   RECT 23.18 695.97 157.32 697.68 ;
   RECT 23.18 697.68 157.32 699.39 ;
   RECT 23.18 699.39 157.32 701.1 ;
   RECT 23.18 701.1 157.32 702.81 ;
   RECT 23.18 702.81 157.32 704.52 ;
   RECT 23.18 704.52 157.32 706.23 ;
   RECT 23.18 706.23 157.32 707.94 ;
   RECT 23.18 707.94 157.32 709.65 ;
   RECT 23.18 709.65 157.32 711.36 ;
   RECT 23.18 711.36 157.32 713.07 ;
   RECT 23.18 713.07 157.32 714.78 ;
   RECT 23.18 714.78 157.32 716.49 ;
   RECT 23.18 716.49 157.32 718.2 ;
   RECT 23.18 718.2 157.32 719.91 ;
   RECT 23.18 719.91 157.32 721.62 ;
   RECT 23.18 721.62 157.32 723.33 ;
   RECT 23.18 723.33 157.32 725.04 ;
   RECT 23.18 725.04 157.32 726.75 ;
   RECT 23.18 726.75 157.32 728.46 ;
   RECT 23.18 728.46 157.32 730.17 ;
   RECT 23.18 730.17 157.32 731.88 ;
   RECT 23.18 731.88 157.32 733.59 ;
   RECT 23.18 733.59 157.32 735.3 ;
   RECT 23.18 735.3 157.32 737.01 ;
   RECT 23.18 737.01 157.32 738.72 ;
   RECT 23.18 738.72 157.32 740.43 ;
   RECT 23.18 740.43 157.32 742.14 ;
   RECT 23.18 742.14 157.32 743.85 ;
   RECT 23.18 743.85 157.32 745.56 ;
   RECT 23.18 745.56 157.32 747.27 ;
   RECT 23.18 747.27 157.32 748.98 ;
   RECT 23.18 748.98 157.32 750.69 ;
   RECT 23.18 750.69 157.32 752.4 ;
   RECT 23.18 752.4 157.32 754.11 ;
 END
END block_414x3969_702

MACRO block_737x819_279
 CLASS BLOCK ;
 FOREIGN block_737x819_279 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 280.06 BY 155.61 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 176.415 153.235 176.985 153.805 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 177.555 153.235 178.125 153.805 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.515 153.235 175.085 153.805 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 170.335 153.235 170.905 153.805 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 171.475 153.235 172.045 153.805 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 168.435 153.235 169.005 153.805 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 145.635 153.235 146.205 153.805 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 144.495 153.235 145.065 153.805 ;
  END
 END o7
 PIN o8
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 139.555 153.235 140.125 153.805 ;
  END
 END o8
 PIN o9
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 138.415 153.235 138.985 153.805 ;
  END
 END o9
 PIN o10
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 151.715 153.235 152.285 153.805 ;
  END
 END o10
 PIN o11
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 150.575 153.235 151.145 153.805 ;
  END
 END o11
 PIN o12
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 148.675 153.235 149.245 153.805 ;
  END
 END o12
 PIN o13
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 269.895 153.235 270.465 153.805 ;
  END
 END o13
 PIN o14
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 271.035 153.235 271.605 153.805 ;
  END
 END o14
 PIN o15
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 267.995 153.235 268.565 153.805 ;
  END
 END o15
 PIN o16
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 263.815 153.235 264.385 153.805 ;
  END
 END o16
 PIN o17
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 264.955 153.235 265.525 153.805 ;
  END
 END o17
 PIN o18
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 261.915 153.235 262.485 153.805 ;
  END
 END o18
 PIN o19
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 257.735 153.235 258.305 153.805 ;
  END
 END o19
 PIN o20
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 258.875 153.235 259.445 153.805 ;
  END
 END o20
 PIN o21
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 255.835 153.235 256.405 153.805 ;
  END
 END o21
 PIN o22
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 251.655 153.235 252.225 153.805 ;
  END
 END o22
 PIN o23
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 252.795 153.235 253.365 153.805 ;
  END
 END o23
 PIN o24
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 249.755 153.235 250.325 153.805 ;
  END
 END o24
 PIN o25
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 245.195 153.235 245.765 153.805 ;
  END
 END o25
 PIN o26
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 247.095 153.235 247.665 153.805 ;
  END
 END o26
 PIN o27
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 244.055 153.235 244.625 153.805 ;
  END
 END o27
 PIN o28
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 233.035 153.235 233.605 153.805 ;
  END
 END o28
 PIN o29
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 231.895 153.235 232.465 153.805 ;
  END
 END o29
 PIN o30
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 229.995 153.235 230.565 153.805 ;
  END
 END o30
 PIN o31
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 226.955 153.235 227.525 153.805 ;
  END
 END o31
 PIN o32
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 225.815 153.235 226.385 153.805 ;
  END
 END o32
 PIN o33
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 242.155 153.235 242.725 153.805 ;
  END
 END o33
 PIN o34
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 237.975 153.235 238.545 153.805 ;
  END
 END o34
 PIN o35
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 239.115 153.235 239.685 153.805 ;
  END
 END o35
 PIN o36
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 236.075 153.235 236.645 153.805 ;
  END
 END o36
 PIN o37
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 162.355 153.235 162.925 153.805 ;
  END
 END o37
 PIN o38
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 136.515 153.235 137.085 153.805 ;
  END
 END o38
 PIN o39
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 223.915 153.235 224.485 153.805 ;
  END
 END o39
 PIN o40
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 180.595 153.235 181.165 153.805 ;
  END
 END o40
 PIN o41
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 156.655 153.235 157.225 153.805 ;
  END
 END o41
 PIN o42
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 182.495 153.235 183.065 153.805 ;
  END
 END o42
 PIN o43
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 164.255 153.235 164.825 153.805 ;
  END
 END o43
 PIN o44
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 241.015 153.235 241.585 153.805 ;
  END
 END o44
 PIN o45
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 179.455 153.235 180.025 153.805 ;
  END
 END o45
 PIN o46
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 165.395 153.235 165.965 153.805 ;
  END
 END o46
 PIN o47
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 266.855 153.235 267.425 153.805 ;
  END
 END o47
 PIN o48
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 260.775 153.235 261.345 153.805 ;
  END
 END o48
 PIN o49
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 254.695 153.235 255.265 153.805 ;
  END
 END o49
 PIN o50
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 185.535 153.235 186.105 153.805 ;
  END
 END o50
 PIN o51
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 159.695 153.235 160.265 153.805 ;
  END
 END o51
 PIN o52
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 173.375 153.235 173.945 153.805 ;
  END
 END o52
 PIN o53
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 234.935 153.235 235.505 153.805 ;
  END
 END o53
 PIN o54
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 141.455 153.235 142.025 153.805 ;
  END
 END o54
 PIN o55
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 167.295 153.235 167.865 153.805 ;
  END
 END o55
 PIN o56
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 228.855 153.235 229.425 153.805 ;
  END
 END o56
 PIN o57
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 153.615 153.235 154.185 153.805 ;
  END
 END o57
 PIN o58
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 142.595 153.235 143.165 153.805 ;
  END
 END o58
 PIN o59
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.755 153.235 155.325 153.805 ;
  END
 END o59
 PIN o60
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 147.535 153.235 148.105 153.805 ;
  END
 END o60
 PIN o61
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 157.795 153.235 158.365 153.805 ;
  END
 END o61
 PIN o62
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 183.635 153.235 184.205 153.805 ;
  END
 END o62
 PIN o63
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 272.935 153.235 273.505 153.805 ;
  END
 END o63
 PIN o64
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 205.295 153.235 205.865 153.805 ;
  END
 END o64
 PIN o65
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.915 0.665 72.485 1.235 ;
  END
 END o65
 PIN o66
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 29.355 153.235 29.925 153.805 ;
  END
 END o66
 PIN o67
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 47.405 3.325 47.975 ;
  END
 END o67
 PIN o68
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 48.165 3.325 48.735 ;
  END
 END o68
 PIN o69
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 103.645 3.325 104.215 ;
  END
 END o69
 PIN o70
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 104.405 3.325 104.975 ;
  END
 END o70
 PIN o71
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 108.015 3.325 108.585 ;
  END
 END o71
 PIN o72
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 108.775 3.325 109.345 ;
  END
 END o72
 PIN o73
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 112.385 3.325 112.955 ;
  END
 END o73
 PIN o74
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 113.145 3.325 113.715 ;
  END
 END o74
 PIN o75
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 116.755 3.325 117.325 ;
  END
 END o75
 PIN o76
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 117.515 3.325 118.085 ;
  END
 END o76
 PIN o77
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 121.125 3.325 121.695 ;
  END
 END o77
 PIN o78
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 121.885 3.325 122.455 ;
  END
 END o78
 PIN o79
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 86.165 3.325 86.735 ;
  END
 END o79
 PIN o80
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 125.495 3.325 126.065 ;
  END
 END o80
 PIN o81
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 126.255 3.325 126.825 ;
  END
 END o81
 PIN o82
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 129.865 3.325 130.435 ;
  END
 END o82
 PIN o83
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 130.625 3.325 131.195 ;
  END
 END o83
 PIN o84
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 134.235 3.325 134.805 ;
  END
 END o84
 PIN o85
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 86.925 3.325 87.495 ;
  END
 END o85
 PIN o86
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 90.535 3.325 91.105 ;
  END
 END o86
 PIN o87
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 91.295 3.325 91.865 ;
  END
 END o87
 PIN o88
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 94.905 3.325 95.475 ;
  END
 END o88
 PIN o89
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 95.665 3.325 96.235 ;
  END
 END o89
 PIN o90
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 99.275 3.325 99.845 ;
  END
 END o90
 PIN o91
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 100.035 3.325 100.605 ;
  END
 END o91
 PIN o92
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 46.835 29.165 47.405 ;
  END
 END o92
 PIN o93
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 49.115 29.165 49.685 ;
  END
 END o93
 PIN o94
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 103.455 29.165 104.025 ;
  END
 END o94
 PIN o95
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 104.785 29.165 105.355 ;
  END
 END o95
 PIN o96
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 107.825 29.165 108.395 ;
  END
 END o96
 PIN o97
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 109.155 29.165 109.725 ;
  END
 END o97
 PIN o98
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 112.195 29.165 112.765 ;
  END
 END o98
 PIN o99
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 113.525 29.165 114.095 ;
  END
 END o99
 PIN o100
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 116.565 29.165 117.135 ;
  END
 END o100
 PIN o101
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 117.895 29.165 118.465 ;
  END
 END o101
 PIN o102
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 120.935 29.165 121.505 ;
  END
 END o102
 PIN o103
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 122.265 29.165 122.835 ;
  END
 END o103
 PIN o104
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 85.975 29.165 86.545 ;
  END
 END o104
 PIN o105
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 125.305 29.165 125.875 ;
  END
 END o105
 PIN o106
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 126.635 29.165 127.205 ;
  END
 END o106
 PIN o107
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 129.675 29.165 130.245 ;
  END
 END o107
 PIN o108
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 131.005 29.165 131.575 ;
  END
 END o108
 PIN o109
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 134.045 29.165 134.615 ;
  END
 END o109
 PIN o110
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 87.305 29.165 87.875 ;
  END
 END o110
 PIN o111
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 90.345 29.165 90.915 ;
  END
 END o111
 PIN o112
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 91.675 29.165 92.245 ;
  END
 END o112
 PIN o113
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 94.715 29.165 95.285 ;
  END
 END o113
 PIN o114
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 96.045 29.165 96.615 ;
  END
 END o114
 PIN o115
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 99.085 29.165 99.655 ;
  END
 END o115
 PIN o116
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 28.595 100.415 29.165 100.985 ;
  END
 END o116
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 44.175 0.665 44.745 1.235 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 43.415 0.665 43.985 1.235 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 54.815 0.665 55.385 1.235 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 42.275 0.665 42.845 1.235 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.575 0.665 56.145 1.235 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 56.335 0.665 56.905 1.235 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 100.795 10.925 101.365 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 98.705 10.925 99.275 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 96.425 10.925 96.995 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 94.335 10.925 94.905 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 92.055 10.925 92.625 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 89.965 10.925 90.535 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 87.685 10.925 88.255 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 85.595 10.925 86.165 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 133.665 10.925 134.235 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 131.385 10.925 131.955 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 127.015 10.925 127.585 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 124.925 10.925 125.495 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 49.115 10.925 49.685 ;
  END
 END i18
 PIN i19
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 122.645 10.925 123.215 ;
  END
 END i19
 PIN i20
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 118.275 10.925 118.845 ;
  END
 END i20
 PIN i21
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 116.185 10.925 116.755 ;
  END
 END i21
 PIN i22
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 113.905 10.925 114.475 ;
  END
 END i22
 PIN i23
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 111.815 10.925 112.385 ;
  END
 END i23
 PIN i24
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 105.165 10.925 105.735 ;
  END
 END i24
 PIN i25
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 103.075 10.925 103.645 ;
  END
 END i25
 PIN i26
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 47.025 10.925 47.595 ;
  END
 END i26
 PIN i27
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 120.555 10.925 121.125 ;
  END
 END i27
 PIN i28
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 129.295 10.925 129.865 ;
  END
 END i28
 PIN i29
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 109.535 10.925 110.105 ;
  END
 END i29
 PIN i30
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 107.445 10.925 108.015 ;
  END
 END i30
 PIN i31
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 59.375 0.665 59.945 1.235 ;
  END
 END i31
 PIN i32
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 37.715 0.665 38.285 1.235 ;
  END
 END i32
 PIN i33
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 35.815 0.665 36.385 1.235 ;
  END
 END i33
 PIN i34
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 60.895 0.665 61.465 1.235 ;
  END
 END i34
 PIN i35
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 39.615 0.665 40.185 1.235 ;
  END
 END i35
 PIN i36
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 34.295 0.665 34.865 1.235 ;
  END
 END i36
 PIN i37
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 70.015 0.665 70.585 1.235 ;
  END
 END i37
 PIN i38
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 0.665 71.725 1.235 ;
  END
 END i38
 PIN i39
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 38.855 0.665 39.425 1.235 ;
  END
 END i39
 PIN i40
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 62.035 0.665 62.605 1.235 ;
  END
 END i40
 PIN i41
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 60.135 0.665 60.705 1.235 ;
  END
 END i41
 PIN i42
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 35.055 0.665 35.625 1.235 ;
  END
 END i42
 PIN i43
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 36.955 0.665 37.525 1.235 ;
  END
 END i43
 PIN i44
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 47.025 4.085 47.595 ;
  END
 END i44
 PIN i45
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 48.735 4.085 49.305 ;
  END
 END i45
 PIN i46
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 103.265 4.085 103.835 ;
  END
 END i46
 PIN i47
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 104.975 4.085 105.545 ;
  END
 END i47
 PIN i48
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 107.635 4.085 108.205 ;
  END
 END i48
 PIN i49
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 109.345 4.085 109.915 ;
  END
 END i49
 PIN i50
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 112.005 4.085 112.575 ;
  END
 END i50
 PIN i51
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 113.715 4.085 114.285 ;
  END
 END i51
 PIN i52
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 116.375 4.085 116.945 ;
  END
 END i52
 PIN i53
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 118.085 4.085 118.655 ;
  END
 END i53
 PIN i54
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 120.745 4.085 121.315 ;
  END
 END i54
 PIN i55
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 122.455 4.085 123.025 ;
  END
 END i55
 PIN i56
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 85.785 4.085 86.355 ;
  END
 END i56
 PIN i57
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 125.115 4.085 125.685 ;
  END
 END i57
 PIN i58
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 126.825 4.085 127.395 ;
  END
 END i58
 PIN i59
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 129.485 4.085 130.055 ;
  END
 END i59
 PIN i60
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 131.195 4.085 131.765 ;
  END
 END i60
 PIN i61
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 133.855 4.085 134.425 ;
  END
 END i61
 PIN i62
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 87.495 4.085 88.065 ;
  END
 END i62
 PIN i63
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 90.155 4.085 90.725 ;
  END
 END i63
 PIN i64
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 91.865 4.085 92.435 ;
  END
 END i64
 PIN i65
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 94.525 4.085 95.095 ;
  END
 END i65
 PIN i66
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 96.235 4.085 96.805 ;
  END
 END i66
 PIN i67
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 98.895 4.085 99.465 ;
  END
 END i67
 PIN i68
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 100.605 4.085 101.175 ;
  END
 END i68
 PIN i69
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 46.455 3.325 47.025 ;
  END
 END i69
 PIN i70
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 49.115 3.325 49.685 ;
  END
 END i70
 PIN i71
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 102.695 3.325 103.265 ;
  END
 END i71
 PIN i72
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 105.355 3.325 105.925 ;
  END
 END i72
 PIN i73
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 107.065 3.325 107.635 ;
  END
 END i73
 PIN i74
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 109.725 3.325 110.295 ;
  END
 END i74
 PIN i75
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 111.435 3.325 112.005 ;
  END
 END i75
 PIN i76
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 114.095 3.325 114.665 ;
  END
 END i76
 PIN i77
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 115.805 3.325 116.375 ;
  END
 END i77
 PIN i78
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 118.465 3.325 119.035 ;
  END
 END i78
 PIN i79
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 120.175 3.325 120.745 ;
  END
 END i79
 PIN i80
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 122.835 3.325 123.405 ;
  END
 END i80
 PIN i81
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 85.215 3.325 85.785 ;
  END
 END i81
 PIN i82
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 124.545 3.325 125.115 ;
  END
 END i82
 PIN i83
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 127.205 3.325 127.775 ;
  END
 END i83
 PIN i84
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 128.915 3.325 129.485 ;
  END
 END i84
 PIN i85
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 131.575 3.325 132.145 ;
  END
 END i85
 PIN i86
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 133.285 3.325 133.855 ;
  END
 END i86
 PIN i87
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 87.875 3.325 88.445 ;
  END
 END i87
 PIN i88
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 89.585 3.325 90.155 ;
  END
 END i88
 PIN i89
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 92.245 3.325 92.815 ;
  END
 END i89
 PIN i90
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 93.955 3.325 94.525 ;
  END
 END i90
 PIN i91
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 96.615 3.325 97.185 ;
  END
 END i91
 PIN i92
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 98.325 3.325 98.895 ;
  END
 END i92
 PIN i93
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 100.985 3.325 101.555 ;
  END
 END i93
 PIN i94
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 65.455 3.325 66.025 ;
  END
 END i94
 PIN i95
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 46.075 4.085 46.645 ;
  END
 END i95
 PIN i96
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 49.685 4.085 50.255 ;
  END
 END i96
 PIN i97
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 102.315 4.085 102.885 ;
  END
 END i97
 PIN i98
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 105.925 4.085 106.495 ;
  END
 END i98
 PIN i99
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 106.685 4.085 107.255 ;
  END
 END i99
 PIN i100
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 110.295 4.085 110.865 ;
  END
 END i100
 PIN i101
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 111.055 4.085 111.625 ;
  END
 END i101
 PIN i102
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 114.665 4.085 115.235 ;
  END
 END i102
 PIN i103
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 115.425 4.085 115.995 ;
  END
 END i103
 PIN i104
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 119.035 4.085 119.605 ;
  END
 END i104
 PIN i105
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 119.795 4.085 120.365 ;
  END
 END i105
 PIN i106
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 123.405 4.085 123.975 ;
  END
 END i106
 PIN i107
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 84.835 4.085 85.405 ;
  END
 END i107
 PIN i108
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 124.165 4.085 124.735 ;
  END
 END i108
 PIN i109
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 127.775 4.085 128.345 ;
  END
 END i109
 PIN i110
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 128.535 4.085 129.105 ;
  END
 END i110
 PIN i111
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 132.145 4.085 132.715 ;
  END
 END i111
 PIN i112
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 132.905 4.085 133.475 ;
  END
 END i112
 PIN i113
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 88.445 4.085 89.015 ;
  END
 END i113
 PIN i114
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 89.205 4.085 89.775 ;
  END
 END i114
 PIN i115
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 92.815 4.085 93.385 ;
  END
 END i115
 PIN i116
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 93.575 4.085 94.145 ;
  END
 END i116
 PIN i117
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 97.185 4.085 97.755 ;
  END
 END i117
 PIN i118
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 97.945 4.085 98.515 ;
  END
 END i118
 PIN i119
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 101.555 4.085 102.125 ;
  END
 END i119
 PIN i120
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 69.255 0.665 69.825 1.235 ;
  END
 END i120
 PIN i121
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 63.935 0.665 64.505 1.235 ;
  END
 END i121
 PIN i122
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 64.695 0.665 65.265 1.235 ;
  END
 END i122
 PIN i123
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 65.455 0.665 66.025 1.235 ;
  END
 END i123
 PIN i124
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 66.595 0.665 67.165 1.235 ;
  END
 END i124
 PIN i125
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 67.355 0.665 67.925 1.235 ;
  END
 END i125
 PIN i126
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 68.495 0.665 69.065 1.235 ;
  END
 END i126
 PIN i127
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 74.575 0.665 75.145 1.235 ;
  END
 END i127
 PIN i128
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 44.935 0.665 45.505 1.235 ;
  END
 END i128
 PIN i129
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 53.675 0.665 54.245 1.235 ;
  END
 END i129
 PIN i130
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 46.075 0.665 46.645 1.235 ;
  END
 END i130
 PIN i131
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 52.915 0.665 53.485 1.235 ;
  END
 END i131
 PIN i132
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 46.835 0.665 47.405 1.235 ;
  END
 END i132
 PIN i133
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 51.775 0.665 52.345 1.235 ;
  END
 END i133
 PIN i134
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 101.175 0.665 101.745 1.235 ;
  END
 END i134
 PIN i135
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 104.595 0.665 105.165 1.235 ;
  END
 END i135
 PIN i136
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 120.175 0.665 120.745 1.235 ;
  END
 END i136
 PIN i137
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 124.735 0.665 125.305 1.235 ;
  END
 END i137
 PIN i138
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 126.635 0.665 127.205 1.235 ;
  END
 END i138
 PIN i139
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 129.295 0.665 129.865 1.235 ;
  END
 END i139
 PIN i140
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 131.195 0.665 131.765 1.235 ;
  END
 END i140
 PIN i141
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 95.855 0.665 96.425 1.235 ;
  END
 END i141
 PIN i142
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 92.815 0.665 93.385 1.235 ;
  END
 END i142
 PIN i143
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 90.155 0.665 90.725 1.235 ;
  END
 END i143
 PIN i144
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 85.595 0.665 86.165 1.235 ;
  END
 END i144
 PIN i145
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 119.415 0.665 119.985 1.235 ;
  END
 END i145
 PIN i146
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 109.155 0.665 109.725 1.235 ;
  END
 END i146
 PIN i147
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 112.955 0.665 113.525 1.235 ;
  END
 END i147
 PIN i148
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 116.755 0.665 117.325 1.235 ;
  END
 END i148
 PIN i149
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 112.195 0.665 112.765 1.235 ;
  END
 END i149
 PIN i150
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 108.395 0.665 108.965 1.235 ;
  END
 END i150
 PIN i151
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 103.835 0.665 104.405 1.235 ;
  END
 END i151
 PIN i152
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 100.035 0.665 100.605 1.235 ;
  END
 END i152
 PIN i153
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 115.615 0.665 116.185 1.235 ;
  END
 END i153
 PIN i154
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 77.995 0.665 78.565 1.235 ;
  END
 END i154
 PIN i155
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 79.135 0.665 79.705 1.235 ;
  END
 END i155
 PIN i156
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 81.795 0.665 82.365 1.235 ;
  END
 END i156
 PIN i157
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 82.935 0.665 83.505 1.235 ;
  END
 END i157
 PIN i158
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 86.355 0.665 86.925 1.235 ;
  END
 END i158
 PIN i159
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 87.495 0.665 88.065 1.235 ;
  END
 END i159
 PIN i160
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 89.015 0.665 89.585 1.235 ;
  END
 END i160
 PIN i161
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 76.095 0.665 76.665 1.235 ;
  END
 END i161
 OBS
  LAYER metal1 ;
   RECT 0 0 280.06 155.61 ;
  LAYER via1 ;
   RECT 0 0 280.06 155.61 ;
  LAYER metal2 ;
   RECT 0 0 280.06 155.61 ;
  LAYER via2 ;
   RECT 0 0 280.06 155.61 ;
  LAYER metal3 ;
   RECT 0 0 280.06 155.61 ;
  LAYER via3 ;
   RECT 0 0 280.06 155.61 ;
  LAYER metal4 ;
   RECT 0 0 280.06 155.61 ;
 END
END block_737x819_279

MACRO block_1100x1557_168
 CLASS BLOCK ;
 FOREIGN block_1100x1557_168 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 418.0 BY 295.83 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 240.825 26.885 241.395 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 248.995 26.885 249.565 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 273.505 26.885 274.075 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 12.635 26.885 13.205 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 20.805 26.885 21.375 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 28.975 26.885 29.545 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 37.145 26.885 37.715 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 45.315 26.885 45.885 ;
  END
 END o7
 PIN o8
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 53.485 26.885 54.055 ;
  END
 END o8
 PIN o9
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 79.895 26.885 80.465 ;
  END
 END o9
 PIN o10
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 281.675 26.885 282.245 ;
  END
 END o10
 PIN o11
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 88.065 26.885 88.635 ;
  END
 END o11
 PIN o12
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 96.235 26.885 96.805 ;
  END
 END o12
 PIN o13
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 104.405 26.885 104.975 ;
  END
 END o13
 PIN o14
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 112.575 26.885 113.145 ;
  END
 END o14
 PIN o15
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 120.745 26.885 121.315 ;
  END
 END o15
 PIN o16
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 128.915 26.885 129.485 ;
  END
 END o16
 PIN o17
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 165.395 26.885 165.965 ;
  END
 END o17
 PIN o18
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 289.845 26.885 290.415 ;
  END
 END o18
 PIN o19
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 257.165 26.885 257.735 ;
  END
 END o19
 PIN o20
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 265.335 26.885 265.905 ;
  END
 END o20
 PIN o21
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 214.415 26.885 214.985 ;
  END
 END o21
 PIN o22
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 181.735 26.885 182.305 ;
  END
 END o22
 PIN o23
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 198.075 26.885 198.645 ;
  END
 END o23
 PIN o24
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 189.905 26.885 190.475 ;
  END
 END o24
 PIN o25
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 206.245 26.885 206.815 ;
  END
 END o25
 PIN o26
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 173.565 26.885 174.135 ;
  END
 END o26
 PIN o27
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 4.465 26.885 5.035 ;
  END
 END o27
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 158.365 3.705 158.935 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 136.705 3.705 137.275 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 141.265 3.705 141.835 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 153.045 3.705 153.615 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 148.675 3.705 149.245 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 157.985 4.465 158.555 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 158.745 4.465 159.315 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 159.125 3.705 159.695 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 149.435 3.705 150.005 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 136.325 4.465 136.895 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 141.645 4.465 142.215 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 144.875 3.705 145.445 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 142.025 3.705 142.595 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 139.935 3.705 140.505 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 137.465 3.705 138.035 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 135.945 3.705 136.515 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 13.015 159.505 13.585 160.075 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 14.535 159.505 15.105 160.075 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 13.015 146.205 13.585 146.775 ;
  END
 END i18
 PIN i19
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 14.535 146.205 15.105 146.775 ;
  END
 END i19
 PIN i20
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 291.555 26.885 292.125 ;
  END
 END i20
 PIN i21
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 283.385 26.885 283.955 ;
  END
 END i21
 PIN i22
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 191.615 26.885 192.185 ;
  END
 END i22
 PIN i23
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 183.445 26.885 184.015 ;
  END
 END i23
 PIN i24
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 175.275 26.885 175.845 ;
  END
 END i24
 PIN i25
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 167.105 26.885 167.675 ;
  END
 END i25
 PIN i26
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 127.205 26.885 127.775 ;
  END
 END i26
 PIN i27
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 119.035 26.885 119.605 ;
  END
 END i27
 PIN i28
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 110.865 26.885 111.435 ;
  END
 END i28
 PIN i29
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 102.695 26.885 103.265 ;
  END
 END i29
 PIN i30
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 94.525 26.885 95.095 ;
  END
 END i30
 PIN i31
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 86.355 26.885 86.925 ;
  END
 END i31
 PIN i32
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 275.215 26.885 275.785 ;
  END
 END i32
 PIN i33
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 78.185 26.885 78.755 ;
  END
 END i33
 PIN i34
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 51.775 26.885 52.345 ;
  END
 END i34
 PIN i35
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 43.605 26.885 44.175 ;
  END
 END i35
 PIN i36
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 35.435 26.885 36.005 ;
  END
 END i36
 PIN i37
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 27.265 26.885 27.835 ;
  END
 END i37
 PIN i38
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 19.095 26.885 19.665 ;
  END
 END i38
 PIN i39
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 10.925 26.885 11.495 ;
  END
 END i39
 PIN i40
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 2.755 26.885 3.325 ;
  END
 END i40
 PIN i41
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 267.045 26.885 267.615 ;
  END
 END i41
 PIN i42
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 258.875 26.885 259.445 ;
  END
 END i42
 PIN i43
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 250.705 26.885 251.275 ;
  END
 END i43
 PIN i44
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 242.535 26.885 243.105 ;
  END
 END i44
 PIN i45
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 216.125 26.885 216.695 ;
  END
 END i45
 PIN i46
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 207.955 26.885 208.525 ;
  END
 END i46
 PIN i47
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 199.785 26.885 200.355 ;
  END
 END i47
 PIN i48
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 260.585 26.885 261.155 ;
  END
 END i48
 PIN i49
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 256.595 27.645 257.165 ;
  END
 END i49
 PIN i50
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 252.415 26.885 252.985 ;
  END
 END i50
 PIN i51
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 268.755 26.885 269.325 ;
  END
 END i51
 PIN i52
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 193.325 26.885 193.895 ;
  END
 END i52
 PIN i53
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 189.335 27.645 189.905 ;
  END
 END i53
 PIN i54
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 185.155 26.885 185.725 ;
  END
 END i54
 PIN i55
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 181.165 27.645 181.735 ;
  END
 END i55
 PIN i56
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 100.985 26.885 101.555 ;
  END
 END i56
 PIN i57
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 104.975 27.645 105.545 ;
  END
 END i57
 PIN i58
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 109.155 26.885 109.725 ;
  END
 END i58
 PIN i59
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 113.145 27.645 113.715 ;
  END
 END i59
 PIN i60
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 33.725 26.885 34.295 ;
  END
 END i60
 PIN i61
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 37.715 27.645 38.285 ;
  END
 END i61
 PIN i62
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 41.895 26.885 42.465 ;
  END
 END i62
 PIN i63
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 25.555 26.885 26.125 ;
  END
 END i63
 PIN i64
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 264.765 27.645 265.335 ;
  END
 END i64
 PIN i65
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 197.505 27.645 198.075 ;
  END
 END i65
 PIN i66
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 96.805 27.645 97.375 ;
  END
 END i66
 PIN i67
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 29.545 27.645 30.115 ;
  END
 END i67
 PIN i68
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 18.335 159.505 18.905 160.075 ;
  END
 END i68
 PIN i69
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 18.335 146.205 18.905 146.775 ;
  END
 END i69
 PIN i70
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 290.985 27.645 291.555 ;
  END
 END i70
 PIN i71
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 282.815 27.645 283.385 ;
  END
 END i71
 PIN i72
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 191.045 27.645 191.615 ;
  END
 END i72
 PIN i73
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 182.875 27.645 183.445 ;
  END
 END i73
 PIN i74
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 174.705 27.645 175.275 ;
  END
 END i74
 PIN i75
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 166.535 27.645 167.105 ;
  END
 END i75
 PIN i76
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 127.775 27.645 128.345 ;
  END
 END i76
 PIN i77
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 119.605 27.645 120.175 ;
  END
 END i77
 PIN i78
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 111.435 27.645 112.005 ;
  END
 END i78
 PIN i79
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 103.265 27.645 103.835 ;
  END
 END i79
 PIN i80
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 95.095 27.645 95.665 ;
  END
 END i80
 PIN i81
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 86.925 27.645 87.495 ;
  END
 END i81
 PIN i82
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 274.645 27.645 275.215 ;
  END
 END i82
 PIN i83
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 78.755 27.645 79.325 ;
  END
 END i83
 PIN i84
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 52.345 27.645 52.915 ;
  END
 END i84
 PIN i85
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 44.175 27.645 44.745 ;
  END
 END i85
 PIN i86
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 36.005 27.645 36.575 ;
  END
 END i86
 PIN i87
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 27.835 27.645 28.405 ;
  END
 END i87
 PIN i88
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 19.665 27.645 20.235 ;
  END
 END i88
 PIN i89
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 11.495 27.645 12.065 ;
  END
 END i89
 PIN i90
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 3.325 27.645 3.895 ;
  END
 END i90
 PIN i91
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 266.475 27.645 267.045 ;
  END
 END i91
 PIN i92
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 258.305 27.645 258.875 ;
  END
 END i92
 PIN i93
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 250.135 27.645 250.705 ;
  END
 END i93
 PIN i94
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 241.965 27.645 242.535 ;
  END
 END i94
 PIN i95
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 215.555 27.645 216.125 ;
  END
 END i95
 PIN i96
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 207.385 27.645 207.955 ;
  END
 END i96
 PIN i97
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 199.215 27.645 199.785 ;
  END
 END i97
 PIN i98
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 151.905 3.705 152.475 ;
  END
 END i98
 PIN i99
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 151.525 4.465 152.095 ;
  END
 END i99
 PIN i100
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 290.415 28.405 290.985 ;
  END
 END i100
 PIN i101
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 282.245 28.405 282.815 ;
  END
 END i101
 PIN i102
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 190.475 28.405 191.045 ;
  END
 END i102
 PIN i103
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 182.305 28.405 182.875 ;
  END
 END i103
 PIN i104
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 174.135 28.405 174.705 ;
  END
 END i104
 PIN i105
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 165.965 28.405 166.535 ;
  END
 END i105
 PIN i106
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 128.345 28.405 128.915 ;
  END
 END i106
 PIN i107
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 120.175 28.405 120.745 ;
  END
 END i107
 PIN i108
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 112.005 28.405 112.575 ;
  END
 END i108
 PIN i109
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 103.835 28.405 104.405 ;
  END
 END i109
 PIN i110
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 95.665 28.405 96.235 ;
  END
 END i110
 PIN i111
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 87.495 28.405 88.065 ;
  END
 END i111
 PIN i112
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 274.075 28.405 274.645 ;
  END
 END i112
 PIN i113
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 79.325 28.405 79.895 ;
  END
 END i113
 PIN i114
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 52.915 28.405 53.485 ;
  END
 END i114
 PIN i115
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 44.745 28.405 45.315 ;
  END
 END i115
 PIN i116
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 36.575 28.405 37.145 ;
  END
 END i116
 PIN i117
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 28.405 28.405 28.975 ;
  END
 END i117
 PIN i118
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 20.235 28.405 20.805 ;
  END
 END i118
 PIN i119
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 12.065 28.405 12.635 ;
  END
 END i119
 PIN i120
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 3.895 28.405 4.465 ;
  END
 END i120
 PIN i121
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 265.905 28.405 266.475 ;
  END
 END i121
 PIN i122
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 257.735 28.405 258.305 ;
  END
 END i122
 PIN i123
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 249.565 28.405 250.135 ;
  END
 END i123
 PIN i124
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 241.395 28.405 241.965 ;
  END
 END i124
 PIN i125
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 214.985 28.405 215.555 ;
  END
 END i125
 PIN i126
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 206.815 28.405 207.385 ;
  END
 END i126
 PIN i127
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 198.645 28.405 199.215 ;
  END
 END i127
 PIN i128
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 4.275 159.505 4.845 160.075 ;
  END
 END i128
 PIN i129
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 5.415 159.505 5.985 160.075 ;
  END
 END i129
 PIN i130
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 7.315 159.505 7.885 160.075 ;
  END
 END i130
 PIN i131
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 8.835 159.505 9.405 160.075 ;
  END
 END i131
 PIN i132
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 159.505 10.925 160.075 ;
  END
 END i132
 PIN i133
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 11.875 159.505 12.445 160.075 ;
  END
 END i133
 PIN i134
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 4.275 146.205 4.845 146.775 ;
  END
 END i134
 PIN i135
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 5.415 146.205 5.985 146.775 ;
  END
 END i135
 PIN i136
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 7.315 146.205 7.885 146.775 ;
  END
 END i136
 PIN i137
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 8.835 146.205 9.405 146.775 ;
  END
 END i137
 PIN i138
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 10.355 146.205 10.925 146.775 ;
  END
 END i138
 PIN i139
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 11.875 146.205 12.445 146.775 ;
  END
 END i139
 OBS
  LAYER metal1 ;
   RECT 23.18 0.0 418.0 1.71 ;
   RECT 23.18 1.71 418.0 3.42 ;
   RECT 23.18 3.42 418.0 5.13 ;
   RECT 23.18 5.13 418.0 6.84 ;
   RECT 23.18 6.84 418.0 8.55 ;
   RECT 23.18 8.55 418.0 10.26 ;
   RECT 23.18 10.26 418.0 11.97 ;
   RECT 23.18 11.97 418.0 13.68 ;
   RECT 23.18 13.68 418.0 15.39 ;
   RECT 23.18 15.39 418.0 17.1 ;
   RECT 23.18 17.1 418.0 18.81 ;
   RECT 23.18 18.81 418.0 20.52 ;
   RECT 23.18 20.52 418.0 22.23 ;
   RECT 23.18 22.23 418.0 23.94 ;
   RECT 23.18 23.94 418.0 25.65 ;
   RECT 23.18 25.65 418.0 27.36 ;
   RECT 23.18 27.36 418.0 29.07 ;
   RECT 23.18 29.07 418.0 30.78 ;
   RECT 23.18 30.78 418.0 32.49 ;
   RECT 23.18 32.49 418.0 34.2 ;
   RECT 23.18 34.2 418.0 35.91 ;
   RECT 23.18 35.91 418.0 37.62 ;
   RECT 23.18 37.62 418.0 39.33 ;
   RECT 23.18 39.33 418.0 41.04 ;
   RECT 23.18 41.04 418.0 42.75 ;
   RECT 23.18 42.75 418.0 44.46 ;
   RECT 23.18 44.46 418.0 46.17 ;
   RECT 23.18 46.17 418.0 47.88 ;
   RECT 23.18 47.88 418.0 49.59 ;
   RECT 23.18 49.59 418.0 51.3 ;
   RECT 23.18 51.3 418.0 53.01 ;
   RECT 23.18 53.01 418.0 54.72 ;
   RECT 23.18 54.72 418.0 56.43 ;
   RECT 23.18 56.43 418.0 58.14 ;
   RECT 23.18 58.14 418.0 59.85 ;
   RECT 23.18 59.85 418.0 61.56 ;
   RECT 23.18 61.56 418.0 63.27 ;
   RECT 23.18 63.27 418.0 64.98 ;
   RECT 23.18 64.98 418.0 66.69 ;
   RECT 23.18 66.69 418.0 68.4 ;
   RECT 23.18 68.4 418.0 70.11 ;
   RECT 23.18 70.11 418.0 71.82 ;
   RECT 23.18 71.82 418.0 73.53 ;
   RECT 23.18 73.53 418.0 75.24 ;
   RECT 23.18 75.24 418.0 76.95 ;
   RECT 23.18 76.95 418.0 78.66 ;
   RECT 23.18 78.66 418.0 80.37 ;
   RECT 23.18 80.37 418.0 82.08 ;
   RECT 23.18 82.08 418.0 83.79 ;
   RECT 23.18 83.79 418.0 85.5 ;
   RECT 23.18 85.5 418.0 87.21 ;
   RECT 23.18 87.21 418.0 88.92 ;
   RECT 23.18 88.92 418.0 90.63 ;
   RECT 23.18 90.63 418.0 92.34 ;
   RECT 23.18 92.34 418.0 94.05 ;
   RECT 23.18 94.05 418.0 95.76 ;
   RECT 23.18 95.76 418.0 97.47 ;
   RECT 23.18 97.47 418.0 99.18 ;
   RECT 23.18 99.18 418.0 100.89 ;
   RECT 23.18 100.89 418.0 102.6 ;
   RECT 23.18 102.6 418.0 104.31 ;
   RECT 23.18 104.31 418.0 106.02 ;
   RECT 23.18 106.02 418.0 107.73 ;
   RECT 23.18 107.73 418.0 109.44 ;
   RECT 23.18 109.44 418.0 111.15 ;
   RECT 23.18 111.15 418.0 112.86 ;
   RECT 23.18 112.86 418.0 114.57 ;
   RECT 23.18 114.57 418.0 116.28 ;
   RECT 23.18 116.28 418.0 117.99 ;
   RECT 23.18 117.99 418.0 119.7 ;
   RECT 23.18 119.7 418.0 121.41 ;
   RECT 23.18 121.41 418.0 123.12 ;
   RECT 23.18 123.12 418.0 124.83 ;
   RECT 23.18 124.83 418.0 126.54 ;
   RECT 23.18 126.54 418.0 128.25 ;
   RECT 23.18 128.25 418.0 129.96 ;
   RECT 23.18 129.96 418.0 131.67 ;
   RECT 23.18 131.67 418.0 133.38 ;
   RECT 0.0 133.38 418.0 135.09 ;
   RECT 0.0 135.09 418.0 136.8 ;
   RECT 0.0 136.8 418.0 138.51 ;
   RECT 0.0 138.51 418.0 140.22 ;
   RECT 0.0 140.22 418.0 141.93 ;
   RECT 0.0 141.93 418.0 143.64 ;
   RECT 0.0 143.64 418.0 145.35 ;
   RECT 0.0 145.35 418.0 147.06 ;
   RECT 0.0 147.06 418.0 148.77 ;
   RECT 0.0 148.77 418.0 150.48 ;
   RECT 0.0 150.48 418.0 152.19 ;
   RECT 0.0 152.19 418.0 153.9 ;
   RECT 0.0 153.9 418.0 155.61 ;
   RECT 0.0 155.61 418.0 157.32 ;
   RECT 0.0 157.32 418.0 159.03 ;
   RECT 0.0 159.03 418.0 160.74 ;
   RECT 0.0 160.74 418.0 162.45 ;
   RECT 23.18 162.45 418.0 164.16 ;
   RECT 23.18 164.16 418.0 165.87 ;
   RECT 23.18 165.87 418.0 167.58 ;
   RECT 23.18 167.58 418.0 169.29 ;
   RECT 23.18 169.29 418.0 171.0 ;
   RECT 23.18 171.0 418.0 172.71 ;
   RECT 23.18 172.71 418.0 174.42 ;
   RECT 23.18 174.42 418.0 176.13 ;
   RECT 23.18 176.13 418.0 177.84 ;
   RECT 23.18 177.84 418.0 179.55 ;
   RECT 23.18 179.55 418.0 181.26 ;
   RECT 23.18 181.26 418.0 182.97 ;
   RECT 23.18 182.97 418.0 184.68 ;
   RECT 23.18 184.68 418.0 186.39 ;
   RECT 23.18 186.39 418.0 188.1 ;
   RECT 23.18 188.1 418.0 189.81 ;
   RECT 23.18 189.81 418.0 191.52 ;
   RECT 23.18 191.52 418.0 193.23 ;
   RECT 23.18 193.23 418.0 194.94 ;
   RECT 23.18 194.94 418.0 196.65 ;
   RECT 23.18 196.65 418.0 198.36 ;
   RECT 23.18 198.36 418.0 200.07 ;
   RECT 23.18 200.07 418.0 201.78 ;
   RECT 23.18 201.78 418.0 203.49 ;
   RECT 23.18 203.49 418.0 205.2 ;
   RECT 23.18 205.2 418.0 206.91 ;
   RECT 23.18 206.91 418.0 208.62 ;
   RECT 23.18 208.62 418.0 210.33 ;
   RECT 23.18 210.33 418.0 212.04 ;
   RECT 23.18 212.04 418.0 213.75 ;
   RECT 23.18 213.75 418.0 215.46 ;
   RECT 23.18 215.46 418.0 217.17 ;
   RECT 23.18 217.17 418.0 218.88 ;
   RECT 23.18 218.88 418.0 220.59 ;
   RECT 23.18 220.59 418.0 222.3 ;
   RECT 23.18 222.3 418.0 224.01 ;
   RECT 23.18 224.01 418.0 225.72 ;
   RECT 23.18 225.72 418.0 227.43 ;
   RECT 23.18 227.43 418.0 229.14 ;
   RECT 23.18 229.14 418.0 230.85 ;
   RECT 23.18 230.85 418.0 232.56 ;
   RECT 23.18 232.56 418.0 234.27 ;
   RECT 23.18 234.27 418.0 235.98 ;
   RECT 23.18 235.98 418.0 237.69 ;
   RECT 23.18 237.69 418.0 239.4 ;
   RECT 23.18 239.4 418.0 241.11 ;
   RECT 23.18 241.11 418.0 242.82 ;
   RECT 23.18 242.82 418.0 244.53 ;
   RECT 23.18 244.53 418.0 246.24 ;
   RECT 23.18 246.24 418.0 247.95 ;
   RECT 23.18 247.95 418.0 249.66 ;
   RECT 23.18 249.66 418.0 251.37 ;
   RECT 23.18 251.37 418.0 253.08 ;
   RECT 23.18 253.08 418.0 254.79 ;
   RECT 23.18 254.79 418.0 256.5 ;
   RECT 23.18 256.5 418.0 258.21 ;
   RECT 23.18 258.21 418.0 259.92 ;
   RECT 23.18 259.92 418.0 261.63 ;
   RECT 23.18 261.63 418.0 263.34 ;
   RECT 23.18 263.34 418.0 265.05 ;
   RECT 23.18 265.05 418.0 266.76 ;
   RECT 23.18 266.76 418.0 268.47 ;
   RECT 23.18 268.47 418.0 270.18 ;
   RECT 23.18 270.18 418.0 271.89 ;
   RECT 23.18 271.89 418.0 273.6 ;
   RECT 23.18 273.6 418.0 275.31 ;
   RECT 23.18 275.31 418.0 277.02 ;
   RECT 23.18 277.02 418.0 278.73 ;
   RECT 23.18 278.73 418.0 280.44 ;
   RECT 23.18 280.44 418.0 282.15 ;
   RECT 23.18 282.15 418.0 283.86 ;
   RECT 23.18 283.86 418.0 285.57 ;
   RECT 23.18 285.57 418.0 287.28 ;
   RECT 23.18 287.28 418.0 288.99 ;
   RECT 23.18 288.99 418.0 290.7 ;
   RECT 23.18 290.7 418.0 292.41 ;
   RECT 23.18 292.41 418.0 294.12 ;
   RECT 23.18 294.12 418.0 295.83 ;
  LAYER via1 ;
   RECT 23.18 0.0 418.0 1.71 ;
   RECT 23.18 1.71 418.0 3.42 ;
   RECT 23.18 3.42 418.0 5.13 ;
   RECT 23.18 5.13 418.0 6.84 ;
   RECT 23.18 6.84 418.0 8.55 ;
   RECT 23.18 8.55 418.0 10.26 ;
   RECT 23.18 10.26 418.0 11.97 ;
   RECT 23.18 11.97 418.0 13.68 ;
   RECT 23.18 13.68 418.0 15.39 ;
   RECT 23.18 15.39 418.0 17.1 ;
   RECT 23.18 17.1 418.0 18.81 ;
   RECT 23.18 18.81 418.0 20.52 ;
   RECT 23.18 20.52 418.0 22.23 ;
   RECT 23.18 22.23 418.0 23.94 ;
   RECT 23.18 23.94 418.0 25.65 ;
   RECT 23.18 25.65 418.0 27.36 ;
   RECT 23.18 27.36 418.0 29.07 ;
   RECT 23.18 29.07 418.0 30.78 ;
   RECT 23.18 30.78 418.0 32.49 ;
   RECT 23.18 32.49 418.0 34.2 ;
   RECT 23.18 34.2 418.0 35.91 ;
   RECT 23.18 35.91 418.0 37.62 ;
   RECT 23.18 37.62 418.0 39.33 ;
   RECT 23.18 39.33 418.0 41.04 ;
   RECT 23.18 41.04 418.0 42.75 ;
   RECT 23.18 42.75 418.0 44.46 ;
   RECT 23.18 44.46 418.0 46.17 ;
   RECT 23.18 46.17 418.0 47.88 ;
   RECT 23.18 47.88 418.0 49.59 ;
   RECT 23.18 49.59 418.0 51.3 ;
   RECT 23.18 51.3 418.0 53.01 ;
   RECT 23.18 53.01 418.0 54.72 ;
   RECT 23.18 54.72 418.0 56.43 ;
   RECT 23.18 56.43 418.0 58.14 ;
   RECT 23.18 58.14 418.0 59.85 ;
   RECT 23.18 59.85 418.0 61.56 ;
   RECT 23.18 61.56 418.0 63.27 ;
   RECT 23.18 63.27 418.0 64.98 ;
   RECT 23.18 64.98 418.0 66.69 ;
   RECT 23.18 66.69 418.0 68.4 ;
   RECT 23.18 68.4 418.0 70.11 ;
   RECT 23.18 70.11 418.0 71.82 ;
   RECT 23.18 71.82 418.0 73.53 ;
   RECT 23.18 73.53 418.0 75.24 ;
   RECT 23.18 75.24 418.0 76.95 ;
   RECT 23.18 76.95 418.0 78.66 ;
   RECT 23.18 78.66 418.0 80.37 ;
   RECT 23.18 80.37 418.0 82.08 ;
   RECT 23.18 82.08 418.0 83.79 ;
   RECT 23.18 83.79 418.0 85.5 ;
   RECT 23.18 85.5 418.0 87.21 ;
   RECT 23.18 87.21 418.0 88.92 ;
   RECT 23.18 88.92 418.0 90.63 ;
   RECT 23.18 90.63 418.0 92.34 ;
   RECT 23.18 92.34 418.0 94.05 ;
   RECT 23.18 94.05 418.0 95.76 ;
   RECT 23.18 95.76 418.0 97.47 ;
   RECT 23.18 97.47 418.0 99.18 ;
   RECT 23.18 99.18 418.0 100.89 ;
   RECT 23.18 100.89 418.0 102.6 ;
   RECT 23.18 102.6 418.0 104.31 ;
   RECT 23.18 104.31 418.0 106.02 ;
   RECT 23.18 106.02 418.0 107.73 ;
   RECT 23.18 107.73 418.0 109.44 ;
   RECT 23.18 109.44 418.0 111.15 ;
   RECT 23.18 111.15 418.0 112.86 ;
   RECT 23.18 112.86 418.0 114.57 ;
   RECT 23.18 114.57 418.0 116.28 ;
   RECT 23.18 116.28 418.0 117.99 ;
   RECT 23.18 117.99 418.0 119.7 ;
   RECT 23.18 119.7 418.0 121.41 ;
   RECT 23.18 121.41 418.0 123.12 ;
   RECT 23.18 123.12 418.0 124.83 ;
   RECT 23.18 124.83 418.0 126.54 ;
   RECT 23.18 126.54 418.0 128.25 ;
   RECT 23.18 128.25 418.0 129.96 ;
   RECT 23.18 129.96 418.0 131.67 ;
   RECT 23.18 131.67 418.0 133.38 ;
   RECT 0.0 133.38 418.0 135.09 ;
   RECT 0.0 135.09 418.0 136.8 ;
   RECT 0.0 136.8 418.0 138.51 ;
   RECT 0.0 138.51 418.0 140.22 ;
   RECT 0.0 140.22 418.0 141.93 ;
   RECT 0.0 141.93 418.0 143.64 ;
   RECT 0.0 143.64 418.0 145.35 ;
   RECT 0.0 145.35 418.0 147.06 ;
   RECT 0.0 147.06 418.0 148.77 ;
   RECT 0.0 148.77 418.0 150.48 ;
   RECT 0.0 150.48 418.0 152.19 ;
   RECT 0.0 152.19 418.0 153.9 ;
   RECT 0.0 153.9 418.0 155.61 ;
   RECT 0.0 155.61 418.0 157.32 ;
   RECT 0.0 157.32 418.0 159.03 ;
   RECT 0.0 159.03 418.0 160.74 ;
   RECT 0.0 160.74 418.0 162.45 ;
   RECT 23.18 162.45 418.0 164.16 ;
   RECT 23.18 164.16 418.0 165.87 ;
   RECT 23.18 165.87 418.0 167.58 ;
   RECT 23.18 167.58 418.0 169.29 ;
   RECT 23.18 169.29 418.0 171.0 ;
   RECT 23.18 171.0 418.0 172.71 ;
   RECT 23.18 172.71 418.0 174.42 ;
   RECT 23.18 174.42 418.0 176.13 ;
   RECT 23.18 176.13 418.0 177.84 ;
   RECT 23.18 177.84 418.0 179.55 ;
   RECT 23.18 179.55 418.0 181.26 ;
   RECT 23.18 181.26 418.0 182.97 ;
   RECT 23.18 182.97 418.0 184.68 ;
   RECT 23.18 184.68 418.0 186.39 ;
   RECT 23.18 186.39 418.0 188.1 ;
   RECT 23.18 188.1 418.0 189.81 ;
   RECT 23.18 189.81 418.0 191.52 ;
   RECT 23.18 191.52 418.0 193.23 ;
   RECT 23.18 193.23 418.0 194.94 ;
   RECT 23.18 194.94 418.0 196.65 ;
   RECT 23.18 196.65 418.0 198.36 ;
   RECT 23.18 198.36 418.0 200.07 ;
   RECT 23.18 200.07 418.0 201.78 ;
   RECT 23.18 201.78 418.0 203.49 ;
   RECT 23.18 203.49 418.0 205.2 ;
   RECT 23.18 205.2 418.0 206.91 ;
   RECT 23.18 206.91 418.0 208.62 ;
   RECT 23.18 208.62 418.0 210.33 ;
   RECT 23.18 210.33 418.0 212.04 ;
   RECT 23.18 212.04 418.0 213.75 ;
   RECT 23.18 213.75 418.0 215.46 ;
   RECT 23.18 215.46 418.0 217.17 ;
   RECT 23.18 217.17 418.0 218.88 ;
   RECT 23.18 218.88 418.0 220.59 ;
   RECT 23.18 220.59 418.0 222.3 ;
   RECT 23.18 222.3 418.0 224.01 ;
   RECT 23.18 224.01 418.0 225.72 ;
   RECT 23.18 225.72 418.0 227.43 ;
   RECT 23.18 227.43 418.0 229.14 ;
   RECT 23.18 229.14 418.0 230.85 ;
   RECT 23.18 230.85 418.0 232.56 ;
   RECT 23.18 232.56 418.0 234.27 ;
   RECT 23.18 234.27 418.0 235.98 ;
   RECT 23.18 235.98 418.0 237.69 ;
   RECT 23.18 237.69 418.0 239.4 ;
   RECT 23.18 239.4 418.0 241.11 ;
   RECT 23.18 241.11 418.0 242.82 ;
   RECT 23.18 242.82 418.0 244.53 ;
   RECT 23.18 244.53 418.0 246.24 ;
   RECT 23.18 246.24 418.0 247.95 ;
   RECT 23.18 247.95 418.0 249.66 ;
   RECT 23.18 249.66 418.0 251.37 ;
   RECT 23.18 251.37 418.0 253.08 ;
   RECT 23.18 253.08 418.0 254.79 ;
   RECT 23.18 254.79 418.0 256.5 ;
   RECT 23.18 256.5 418.0 258.21 ;
   RECT 23.18 258.21 418.0 259.92 ;
   RECT 23.18 259.92 418.0 261.63 ;
   RECT 23.18 261.63 418.0 263.34 ;
   RECT 23.18 263.34 418.0 265.05 ;
   RECT 23.18 265.05 418.0 266.76 ;
   RECT 23.18 266.76 418.0 268.47 ;
   RECT 23.18 268.47 418.0 270.18 ;
   RECT 23.18 270.18 418.0 271.89 ;
   RECT 23.18 271.89 418.0 273.6 ;
   RECT 23.18 273.6 418.0 275.31 ;
   RECT 23.18 275.31 418.0 277.02 ;
   RECT 23.18 277.02 418.0 278.73 ;
   RECT 23.18 278.73 418.0 280.44 ;
   RECT 23.18 280.44 418.0 282.15 ;
   RECT 23.18 282.15 418.0 283.86 ;
   RECT 23.18 283.86 418.0 285.57 ;
   RECT 23.18 285.57 418.0 287.28 ;
   RECT 23.18 287.28 418.0 288.99 ;
   RECT 23.18 288.99 418.0 290.7 ;
   RECT 23.18 290.7 418.0 292.41 ;
   RECT 23.18 292.41 418.0 294.12 ;
   RECT 23.18 294.12 418.0 295.83 ;
  LAYER metal2 ;
   RECT 23.18 0.0 418.0 1.71 ;
   RECT 23.18 1.71 418.0 3.42 ;
   RECT 23.18 3.42 418.0 5.13 ;
   RECT 23.18 5.13 418.0 6.84 ;
   RECT 23.18 6.84 418.0 8.55 ;
   RECT 23.18 8.55 418.0 10.26 ;
   RECT 23.18 10.26 418.0 11.97 ;
   RECT 23.18 11.97 418.0 13.68 ;
   RECT 23.18 13.68 418.0 15.39 ;
   RECT 23.18 15.39 418.0 17.1 ;
   RECT 23.18 17.1 418.0 18.81 ;
   RECT 23.18 18.81 418.0 20.52 ;
   RECT 23.18 20.52 418.0 22.23 ;
   RECT 23.18 22.23 418.0 23.94 ;
   RECT 23.18 23.94 418.0 25.65 ;
   RECT 23.18 25.65 418.0 27.36 ;
   RECT 23.18 27.36 418.0 29.07 ;
   RECT 23.18 29.07 418.0 30.78 ;
   RECT 23.18 30.78 418.0 32.49 ;
   RECT 23.18 32.49 418.0 34.2 ;
   RECT 23.18 34.2 418.0 35.91 ;
   RECT 23.18 35.91 418.0 37.62 ;
   RECT 23.18 37.62 418.0 39.33 ;
   RECT 23.18 39.33 418.0 41.04 ;
   RECT 23.18 41.04 418.0 42.75 ;
   RECT 23.18 42.75 418.0 44.46 ;
   RECT 23.18 44.46 418.0 46.17 ;
   RECT 23.18 46.17 418.0 47.88 ;
   RECT 23.18 47.88 418.0 49.59 ;
   RECT 23.18 49.59 418.0 51.3 ;
   RECT 23.18 51.3 418.0 53.01 ;
   RECT 23.18 53.01 418.0 54.72 ;
   RECT 23.18 54.72 418.0 56.43 ;
   RECT 23.18 56.43 418.0 58.14 ;
   RECT 23.18 58.14 418.0 59.85 ;
   RECT 23.18 59.85 418.0 61.56 ;
   RECT 23.18 61.56 418.0 63.27 ;
   RECT 23.18 63.27 418.0 64.98 ;
   RECT 23.18 64.98 418.0 66.69 ;
   RECT 23.18 66.69 418.0 68.4 ;
   RECT 23.18 68.4 418.0 70.11 ;
   RECT 23.18 70.11 418.0 71.82 ;
   RECT 23.18 71.82 418.0 73.53 ;
   RECT 23.18 73.53 418.0 75.24 ;
   RECT 23.18 75.24 418.0 76.95 ;
   RECT 23.18 76.95 418.0 78.66 ;
   RECT 23.18 78.66 418.0 80.37 ;
   RECT 23.18 80.37 418.0 82.08 ;
   RECT 23.18 82.08 418.0 83.79 ;
   RECT 23.18 83.79 418.0 85.5 ;
   RECT 23.18 85.5 418.0 87.21 ;
   RECT 23.18 87.21 418.0 88.92 ;
   RECT 23.18 88.92 418.0 90.63 ;
   RECT 23.18 90.63 418.0 92.34 ;
   RECT 23.18 92.34 418.0 94.05 ;
   RECT 23.18 94.05 418.0 95.76 ;
   RECT 23.18 95.76 418.0 97.47 ;
   RECT 23.18 97.47 418.0 99.18 ;
   RECT 23.18 99.18 418.0 100.89 ;
   RECT 23.18 100.89 418.0 102.6 ;
   RECT 23.18 102.6 418.0 104.31 ;
   RECT 23.18 104.31 418.0 106.02 ;
   RECT 23.18 106.02 418.0 107.73 ;
   RECT 23.18 107.73 418.0 109.44 ;
   RECT 23.18 109.44 418.0 111.15 ;
   RECT 23.18 111.15 418.0 112.86 ;
   RECT 23.18 112.86 418.0 114.57 ;
   RECT 23.18 114.57 418.0 116.28 ;
   RECT 23.18 116.28 418.0 117.99 ;
   RECT 23.18 117.99 418.0 119.7 ;
   RECT 23.18 119.7 418.0 121.41 ;
   RECT 23.18 121.41 418.0 123.12 ;
   RECT 23.18 123.12 418.0 124.83 ;
   RECT 23.18 124.83 418.0 126.54 ;
   RECT 23.18 126.54 418.0 128.25 ;
   RECT 23.18 128.25 418.0 129.96 ;
   RECT 23.18 129.96 418.0 131.67 ;
   RECT 23.18 131.67 418.0 133.38 ;
   RECT 0.0 133.38 418.0 135.09 ;
   RECT 0.0 135.09 418.0 136.8 ;
   RECT 0.0 136.8 418.0 138.51 ;
   RECT 0.0 138.51 418.0 140.22 ;
   RECT 0.0 140.22 418.0 141.93 ;
   RECT 0.0 141.93 418.0 143.64 ;
   RECT 0.0 143.64 418.0 145.35 ;
   RECT 0.0 145.35 418.0 147.06 ;
   RECT 0.0 147.06 418.0 148.77 ;
   RECT 0.0 148.77 418.0 150.48 ;
   RECT 0.0 150.48 418.0 152.19 ;
   RECT 0.0 152.19 418.0 153.9 ;
   RECT 0.0 153.9 418.0 155.61 ;
   RECT 0.0 155.61 418.0 157.32 ;
   RECT 0.0 157.32 418.0 159.03 ;
   RECT 0.0 159.03 418.0 160.74 ;
   RECT 0.0 160.74 418.0 162.45 ;
   RECT 23.18 162.45 418.0 164.16 ;
   RECT 23.18 164.16 418.0 165.87 ;
   RECT 23.18 165.87 418.0 167.58 ;
   RECT 23.18 167.58 418.0 169.29 ;
   RECT 23.18 169.29 418.0 171.0 ;
   RECT 23.18 171.0 418.0 172.71 ;
   RECT 23.18 172.71 418.0 174.42 ;
   RECT 23.18 174.42 418.0 176.13 ;
   RECT 23.18 176.13 418.0 177.84 ;
   RECT 23.18 177.84 418.0 179.55 ;
   RECT 23.18 179.55 418.0 181.26 ;
   RECT 23.18 181.26 418.0 182.97 ;
   RECT 23.18 182.97 418.0 184.68 ;
   RECT 23.18 184.68 418.0 186.39 ;
   RECT 23.18 186.39 418.0 188.1 ;
   RECT 23.18 188.1 418.0 189.81 ;
   RECT 23.18 189.81 418.0 191.52 ;
   RECT 23.18 191.52 418.0 193.23 ;
   RECT 23.18 193.23 418.0 194.94 ;
   RECT 23.18 194.94 418.0 196.65 ;
   RECT 23.18 196.65 418.0 198.36 ;
   RECT 23.18 198.36 418.0 200.07 ;
   RECT 23.18 200.07 418.0 201.78 ;
   RECT 23.18 201.78 418.0 203.49 ;
   RECT 23.18 203.49 418.0 205.2 ;
   RECT 23.18 205.2 418.0 206.91 ;
   RECT 23.18 206.91 418.0 208.62 ;
   RECT 23.18 208.62 418.0 210.33 ;
   RECT 23.18 210.33 418.0 212.04 ;
   RECT 23.18 212.04 418.0 213.75 ;
   RECT 23.18 213.75 418.0 215.46 ;
   RECT 23.18 215.46 418.0 217.17 ;
   RECT 23.18 217.17 418.0 218.88 ;
   RECT 23.18 218.88 418.0 220.59 ;
   RECT 23.18 220.59 418.0 222.3 ;
   RECT 23.18 222.3 418.0 224.01 ;
   RECT 23.18 224.01 418.0 225.72 ;
   RECT 23.18 225.72 418.0 227.43 ;
   RECT 23.18 227.43 418.0 229.14 ;
   RECT 23.18 229.14 418.0 230.85 ;
   RECT 23.18 230.85 418.0 232.56 ;
   RECT 23.18 232.56 418.0 234.27 ;
   RECT 23.18 234.27 418.0 235.98 ;
   RECT 23.18 235.98 418.0 237.69 ;
   RECT 23.18 237.69 418.0 239.4 ;
   RECT 23.18 239.4 418.0 241.11 ;
   RECT 23.18 241.11 418.0 242.82 ;
   RECT 23.18 242.82 418.0 244.53 ;
   RECT 23.18 244.53 418.0 246.24 ;
   RECT 23.18 246.24 418.0 247.95 ;
   RECT 23.18 247.95 418.0 249.66 ;
   RECT 23.18 249.66 418.0 251.37 ;
   RECT 23.18 251.37 418.0 253.08 ;
   RECT 23.18 253.08 418.0 254.79 ;
   RECT 23.18 254.79 418.0 256.5 ;
   RECT 23.18 256.5 418.0 258.21 ;
   RECT 23.18 258.21 418.0 259.92 ;
   RECT 23.18 259.92 418.0 261.63 ;
   RECT 23.18 261.63 418.0 263.34 ;
   RECT 23.18 263.34 418.0 265.05 ;
   RECT 23.18 265.05 418.0 266.76 ;
   RECT 23.18 266.76 418.0 268.47 ;
   RECT 23.18 268.47 418.0 270.18 ;
   RECT 23.18 270.18 418.0 271.89 ;
   RECT 23.18 271.89 418.0 273.6 ;
   RECT 23.18 273.6 418.0 275.31 ;
   RECT 23.18 275.31 418.0 277.02 ;
   RECT 23.18 277.02 418.0 278.73 ;
   RECT 23.18 278.73 418.0 280.44 ;
   RECT 23.18 280.44 418.0 282.15 ;
   RECT 23.18 282.15 418.0 283.86 ;
   RECT 23.18 283.86 418.0 285.57 ;
   RECT 23.18 285.57 418.0 287.28 ;
   RECT 23.18 287.28 418.0 288.99 ;
   RECT 23.18 288.99 418.0 290.7 ;
   RECT 23.18 290.7 418.0 292.41 ;
   RECT 23.18 292.41 418.0 294.12 ;
   RECT 23.18 294.12 418.0 295.83 ;
  LAYER via2 ;
   RECT 23.18 0.0 418.0 1.71 ;
   RECT 23.18 1.71 418.0 3.42 ;
   RECT 23.18 3.42 418.0 5.13 ;
   RECT 23.18 5.13 418.0 6.84 ;
   RECT 23.18 6.84 418.0 8.55 ;
   RECT 23.18 8.55 418.0 10.26 ;
   RECT 23.18 10.26 418.0 11.97 ;
   RECT 23.18 11.97 418.0 13.68 ;
   RECT 23.18 13.68 418.0 15.39 ;
   RECT 23.18 15.39 418.0 17.1 ;
   RECT 23.18 17.1 418.0 18.81 ;
   RECT 23.18 18.81 418.0 20.52 ;
   RECT 23.18 20.52 418.0 22.23 ;
   RECT 23.18 22.23 418.0 23.94 ;
   RECT 23.18 23.94 418.0 25.65 ;
   RECT 23.18 25.65 418.0 27.36 ;
   RECT 23.18 27.36 418.0 29.07 ;
   RECT 23.18 29.07 418.0 30.78 ;
   RECT 23.18 30.78 418.0 32.49 ;
   RECT 23.18 32.49 418.0 34.2 ;
   RECT 23.18 34.2 418.0 35.91 ;
   RECT 23.18 35.91 418.0 37.62 ;
   RECT 23.18 37.62 418.0 39.33 ;
   RECT 23.18 39.33 418.0 41.04 ;
   RECT 23.18 41.04 418.0 42.75 ;
   RECT 23.18 42.75 418.0 44.46 ;
   RECT 23.18 44.46 418.0 46.17 ;
   RECT 23.18 46.17 418.0 47.88 ;
   RECT 23.18 47.88 418.0 49.59 ;
   RECT 23.18 49.59 418.0 51.3 ;
   RECT 23.18 51.3 418.0 53.01 ;
   RECT 23.18 53.01 418.0 54.72 ;
   RECT 23.18 54.72 418.0 56.43 ;
   RECT 23.18 56.43 418.0 58.14 ;
   RECT 23.18 58.14 418.0 59.85 ;
   RECT 23.18 59.85 418.0 61.56 ;
   RECT 23.18 61.56 418.0 63.27 ;
   RECT 23.18 63.27 418.0 64.98 ;
   RECT 23.18 64.98 418.0 66.69 ;
   RECT 23.18 66.69 418.0 68.4 ;
   RECT 23.18 68.4 418.0 70.11 ;
   RECT 23.18 70.11 418.0 71.82 ;
   RECT 23.18 71.82 418.0 73.53 ;
   RECT 23.18 73.53 418.0 75.24 ;
   RECT 23.18 75.24 418.0 76.95 ;
   RECT 23.18 76.95 418.0 78.66 ;
   RECT 23.18 78.66 418.0 80.37 ;
   RECT 23.18 80.37 418.0 82.08 ;
   RECT 23.18 82.08 418.0 83.79 ;
   RECT 23.18 83.79 418.0 85.5 ;
   RECT 23.18 85.5 418.0 87.21 ;
   RECT 23.18 87.21 418.0 88.92 ;
   RECT 23.18 88.92 418.0 90.63 ;
   RECT 23.18 90.63 418.0 92.34 ;
   RECT 23.18 92.34 418.0 94.05 ;
   RECT 23.18 94.05 418.0 95.76 ;
   RECT 23.18 95.76 418.0 97.47 ;
   RECT 23.18 97.47 418.0 99.18 ;
   RECT 23.18 99.18 418.0 100.89 ;
   RECT 23.18 100.89 418.0 102.6 ;
   RECT 23.18 102.6 418.0 104.31 ;
   RECT 23.18 104.31 418.0 106.02 ;
   RECT 23.18 106.02 418.0 107.73 ;
   RECT 23.18 107.73 418.0 109.44 ;
   RECT 23.18 109.44 418.0 111.15 ;
   RECT 23.18 111.15 418.0 112.86 ;
   RECT 23.18 112.86 418.0 114.57 ;
   RECT 23.18 114.57 418.0 116.28 ;
   RECT 23.18 116.28 418.0 117.99 ;
   RECT 23.18 117.99 418.0 119.7 ;
   RECT 23.18 119.7 418.0 121.41 ;
   RECT 23.18 121.41 418.0 123.12 ;
   RECT 23.18 123.12 418.0 124.83 ;
   RECT 23.18 124.83 418.0 126.54 ;
   RECT 23.18 126.54 418.0 128.25 ;
   RECT 23.18 128.25 418.0 129.96 ;
   RECT 23.18 129.96 418.0 131.67 ;
   RECT 23.18 131.67 418.0 133.38 ;
   RECT 0.0 133.38 418.0 135.09 ;
   RECT 0.0 135.09 418.0 136.8 ;
   RECT 0.0 136.8 418.0 138.51 ;
   RECT 0.0 138.51 418.0 140.22 ;
   RECT 0.0 140.22 418.0 141.93 ;
   RECT 0.0 141.93 418.0 143.64 ;
   RECT 0.0 143.64 418.0 145.35 ;
   RECT 0.0 145.35 418.0 147.06 ;
   RECT 0.0 147.06 418.0 148.77 ;
   RECT 0.0 148.77 418.0 150.48 ;
   RECT 0.0 150.48 418.0 152.19 ;
   RECT 0.0 152.19 418.0 153.9 ;
   RECT 0.0 153.9 418.0 155.61 ;
   RECT 0.0 155.61 418.0 157.32 ;
   RECT 0.0 157.32 418.0 159.03 ;
   RECT 0.0 159.03 418.0 160.74 ;
   RECT 0.0 160.74 418.0 162.45 ;
   RECT 23.18 162.45 418.0 164.16 ;
   RECT 23.18 164.16 418.0 165.87 ;
   RECT 23.18 165.87 418.0 167.58 ;
   RECT 23.18 167.58 418.0 169.29 ;
   RECT 23.18 169.29 418.0 171.0 ;
   RECT 23.18 171.0 418.0 172.71 ;
   RECT 23.18 172.71 418.0 174.42 ;
   RECT 23.18 174.42 418.0 176.13 ;
   RECT 23.18 176.13 418.0 177.84 ;
   RECT 23.18 177.84 418.0 179.55 ;
   RECT 23.18 179.55 418.0 181.26 ;
   RECT 23.18 181.26 418.0 182.97 ;
   RECT 23.18 182.97 418.0 184.68 ;
   RECT 23.18 184.68 418.0 186.39 ;
   RECT 23.18 186.39 418.0 188.1 ;
   RECT 23.18 188.1 418.0 189.81 ;
   RECT 23.18 189.81 418.0 191.52 ;
   RECT 23.18 191.52 418.0 193.23 ;
   RECT 23.18 193.23 418.0 194.94 ;
   RECT 23.18 194.94 418.0 196.65 ;
   RECT 23.18 196.65 418.0 198.36 ;
   RECT 23.18 198.36 418.0 200.07 ;
   RECT 23.18 200.07 418.0 201.78 ;
   RECT 23.18 201.78 418.0 203.49 ;
   RECT 23.18 203.49 418.0 205.2 ;
   RECT 23.18 205.2 418.0 206.91 ;
   RECT 23.18 206.91 418.0 208.62 ;
   RECT 23.18 208.62 418.0 210.33 ;
   RECT 23.18 210.33 418.0 212.04 ;
   RECT 23.18 212.04 418.0 213.75 ;
   RECT 23.18 213.75 418.0 215.46 ;
   RECT 23.18 215.46 418.0 217.17 ;
   RECT 23.18 217.17 418.0 218.88 ;
   RECT 23.18 218.88 418.0 220.59 ;
   RECT 23.18 220.59 418.0 222.3 ;
   RECT 23.18 222.3 418.0 224.01 ;
   RECT 23.18 224.01 418.0 225.72 ;
   RECT 23.18 225.72 418.0 227.43 ;
   RECT 23.18 227.43 418.0 229.14 ;
   RECT 23.18 229.14 418.0 230.85 ;
   RECT 23.18 230.85 418.0 232.56 ;
   RECT 23.18 232.56 418.0 234.27 ;
   RECT 23.18 234.27 418.0 235.98 ;
   RECT 23.18 235.98 418.0 237.69 ;
   RECT 23.18 237.69 418.0 239.4 ;
   RECT 23.18 239.4 418.0 241.11 ;
   RECT 23.18 241.11 418.0 242.82 ;
   RECT 23.18 242.82 418.0 244.53 ;
   RECT 23.18 244.53 418.0 246.24 ;
   RECT 23.18 246.24 418.0 247.95 ;
   RECT 23.18 247.95 418.0 249.66 ;
   RECT 23.18 249.66 418.0 251.37 ;
   RECT 23.18 251.37 418.0 253.08 ;
   RECT 23.18 253.08 418.0 254.79 ;
   RECT 23.18 254.79 418.0 256.5 ;
   RECT 23.18 256.5 418.0 258.21 ;
   RECT 23.18 258.21 418.0 259.92 ;
   RECT 23.18 259.92 418.0 261.63 ;
   RECT 23.18 261.63 418.0 263.34 ;
   RECT 23.18 263.34 418.0 265.05 ;
   RECT 23.18 265.05 418.0 266.76 ;
   RECT 23.18 266.76 418.0 268.47 ;
   RECT 23.18 268.47 418.0 270.18 ;
   RECT 23.18 270.18 418.0 271.89 ;
   RECT 23.18 271.89 418.0 273.6 ;
   RECT 23.18 273.6 418.0 275.31 ;
   RECT 23.18 275.31 418.0 277.02 ;
   RECT 23.18 277.02 418.0 278.73 ;
   RECT 23.18 278.73 418.0 280.44 ;
   RECT 23.18 280.44 418.0 282.15 ;
   RECT 23.18 282.15 418.0 283.86 ;
   RECT 23.18 283.86 418.0 285.57 ;
   RECT 23.18 285.57 418.0 287.28 ;
   RECT 23.18 287.28 418.0 288.99 ;
   RECT 23.18 288.99 418.0 290.7 ;
   RECT 23.18 290.7 418.0 292.41 ;
   RECT 23.18 292.41 418.0 294.12 ;
   RECT 23.18 294.12 418.0 295.83 ;
  LAYER metal3 ;
   RECT 23.18 0.0 418.0 1.71 ;
   RECT 23.18 1.71 418.0 3.42 ;
   RECT 23.18 3.42 418.0 5.13 ;
   RECT 23.18 5.13 418.0 6.84 ;
   RECT 23.18 6.84 418.0 8.55 ;
   RECT 23.18 8.55 418.0 10.26 ;
   RECT 23.18 10.26 418.0 11.97 ;
   RECT 23.18 11.97 418.0 13.68 ;
   RECT 23.18 13.68 418.0 15.39 ;
   RECT 23.18 15.39 418.0 17.1 ;
   RECT 23.18 17.1 418.0 18.81 ;
   RECT 23.18 18.81 418.0 20.52 ;
   RECT 23.18 20.52 418.0 22.23 ;
   RECT 23.18 22.23 418.0 23.94 ;
   RECT 23.18 23.94 418.0 25.65 ;
   RECT 23.18 25.65 418.0 27.36 ;
   RECT 23.18 27.36 418.0 29.07 ;
   RECT 23.18 29.07 418.0 30.78 ;
   RECT 23.18 30.78 418.0 32.49 ;
   RECT 23.18 32.49 418.0 34.2 ;
   RECT 23.18 34.2 418.0 35.91 ;
   RECT 23.18 35.91 418.0 37.62 ;
   RECT 23.18 37.62 418.0 39.33 ;
   RECT 23.18 39.33 418.0 41.04 ;
   RECT 23.18 41.04 418.0 42.75 ;
   RECT 23.18 42.75 418.0 44.46 ;
   RECT 23.18 44.46 418.0 46.17 ;
   RECT 23.18 46.17 418.0 47.88 ;
   RECT 23.18 47.88 418.0 49.59 ;
   RECT 23.18 49.59 418.0 51.3 ;
   RECT 23.18 51.3 418.0 53.01 ;
   RECT 23.18 53.01 418.0 54.72 ;
   RECT 23.18 54.72 418.0 56.43 ;
   RECT 23.18 56.43 418.0 58.14 ;
   RECT 23.18 58.14 418.0 59.85 ;
   RECT 23.18 59.85 418.0 61.56 ;
   RECT 23.18 61.56 418.0 63.27 ;
   RECT 23.18 63.27 418.0 64.98 ;
   RECT 23.18 64.98 418.0 66.69 ;
   RECT 23.18 66.69 418.0 68.4 ;
   RECT 23.18 68.4 418.0 70.11 ;
   RECT 23.18 70.11 418.0 71.82 ;
   RECT 23.18 71.82 418.0 73.53 ;
   RECT 23.18 73.53 418.0 75.24 ;
   RECT 23.18 75.24 418.0 76.95 ;
   RECT 23.18 76.95 418.0 78.66 ;
   RECT 23.18 78.66 418.0 80.37 ;
   RECT 23.18 80.37 418.0 82.08 ;
   RECT 23.18 82.08 418.0 83.79 ;
   RECT 23.18 83.79 418.0 85.5 ;
   RECT 23.18 85.5 418.0 87.21 ;
   RECT 23.18 87.21 418.0 88.92 ;
   RECT 23.18 88.92 418.0 90.63 ;
   RECT 23.18 90.63 418.0 92.34 ;
   RECT 23.18 92.34 418.0 94.05 ;
   RECT 23.18 94.05 418.0 95.76 ;
   RECT 23.18 95.76 418.0 97.47 ;
   RECT 23.18 97.47 418.0 99.18 ;
   RECT 23.18 99.18 418.0 100.89 ;
   RECT 23.18 100.89 418.0 102.6 ;
   RECT 23.18 102.6 418.0 104.31 ;
   RECT 23.18 104.31 418.0 106.02 ;
   RECT 23.18 106.02 418.0 107.73 ;
   RECT 23.18 107.73 418.0 109.44 ;
   RECT 23.18 109.44 418.0 111.15 ;
   RECT 23.18 111.15 418.0 112.86 ;
   RECT 23.18 112.86 418.0 114.57 ;
   RECT 23.18 114.57 418.0 116.28 ;
   RECT 23.18 116.28 418.0 117.99 ;
   RECT 23.18 117.99 418.0 119.7 ;
   RECT 23.18 119.7 418.0 121.41 ;
   RECT 23.18 121.41 418.0 123.12 ;
   RECT 23.18 123.12 418.0 124.83 ;
   RECT 23.18 124.83 418.0 126.54 ;
   RECT 23.18 126.54 418.0 128.25 ;
   RECT 23.18 128.25 418.0 129.96 ;
   RECT 23.18 129.96 418.0 131.67 ;
   RECT 23.18 131.67 418.0 133.38 ;
   RECT 0.0 133.38 418.0 135.09 ;
   RECT 0.0 135.09 418.0 136.8 ;
   RECT 0.0 136.8 418.0 138.51 ;
   RECT 0.0 138.51 418.0 140.22 ;
   RECT 0.0 140.22 418.0 141.93 ;
   RECT 0.0 141.93 418.0 143.64 ;
   RECT 0.0 143.64 418.0 145.35 ;
   RECT 0.0 145.35 418.0 147.06 ;
   RECT 0.0 147.06 418.0 148.77 ;
   RECT 0.0 148.77 418.0 150.48 ;
   RECT 0.0 150.48 418.0 152.19 ;
   RECT 0.0 152.19 418.0 153.9 ;
   RECT 0.0 153.9 418.0 155.61 ;
   RECT 0.0 155.61 418.0 157.32 ;
   RECT 0.0 157.32 418.0 159.03 ;
   RECT 0.0 159.03 418.0 160.74 ;
   RECT 0.0 160.74 418.0 162.45 ;
   RECT 23.18 162.45 418.0 164.16 ;
   RECT 23.18 164.16 418.0 165.87 ;
   RECT 23.18 165.87 418.0 167.58 ;
   RECT 23.18 167.58 418.0 169.29 ;
   RECT 23.18 169.29 418.0 171.0 ;
   RECT 23.18 171.0 418.0 172.71 ;
   RECT 23.18 172.71 418.0 174.42 ;
   RECT 23.18 174.42 418.0 176.13 ;
   RECT 23.18 176.13 418.0 177.84 ;
   RECT 23.18 177.84 418.0 179.55 ;
   RECT 23.18 179.55 418.0 181.26 ;
   RECT 23.18 181.26 418.0 182.97 ;
   RECT 23.18 182.97 418.0 184.68 ;
   RECT 23.18 184.68 418.0 186.39 ;
   RECT 23.18 186.39 418.0 188.1 ;
   RECT 23.18 188.1 418.0 189.81 ;
   RECT 23.18 189.81 418.0 191.52 ;
   RECT 23.18 191.52 418.0 193.23 ;
   RECT 23.18 193.23 418.0 194.94 ;
   RECT 23.18 194.94 418.0 196.65 ;
   RECT 23.18 196.65 418.0 198.36 ;
   RECT 23.18 198.36 418.0 200.07 ;
   RECT 23.18 200.07 418.0 201.78 ;
   RECT 23.18 201.78 418.0 203.49 ;
   RECT 23.18 203.49 418.0 205.2 ;
   RECT 23.18 205.2 418.0 206.91 ;
   RECT 23.18 206.91 418.0 208.62 ;
   RECT 23.18 208.62 418.0 210.33 ;
   RECT 23.18 210.33 418.0 212.04 ;
   RECT 23.18 212.04 418.0 213.75 ;
   RECT 23.18 213.75 418.0 215.46 ;
   RECT 23.18 215.46 418.0 217.17 ;
   RECT 23.18 217.17 418.0 218.88 ;
   RECT 23.18 218.88 418.0 220.59 ;
   RECT 23.18 220.59 418.0 222.3 ;
   RECT 23.18 222.3 418.0 224.01 ;
   RECT 23.18 224.01 418.0 225.72 ;
   RECT 23.18 225.72 418.0 227.43 ;
   RECT 23.18 227.43 418.0 229.14 ;
   RECT 23.18 229.14 418.0 230.85 ;
   RECT 23.18 230.85 418.0 232.56 ;
   RECT 23.18 232.56 418.0 234.27 ;
   RECT 23.18 234.27 418.0 235.98 ;
   RECT 23.18 235.98 418.0 237.69 ;
   RECT 23.18 237.69 418.0 239.4 ;
   RECT 23.18 239.4 418.0 241.11 ;
   RECT 23.18 241.11 418.0 242.82 ;
   RECT 23.18 242.82 418.0 244.53 ;
   RECT 23.18 244.53 418.0 246.24 ;
   RECT 23.18 246.24 418.0 247.95 ;
   RECT 23.18 247.95 418.0 249.66 ;
   RECT 23.18 249.66 418.0 251.37 ;
   RECT 23.18 251.37 418.0 253.08 ;
   RECT 23.18 253.08 418.0 254.79 ;
   RECT 23.18 254.79 418.0 256.5 ;
   RECT 23.18 256.5 418.0 258.21 ;
   RECT 23.18 258.21 418.0 259.92 ;
   RECT 23.18 259.92 418.0 261.63 ;
   RECT 23.18 261.63 418.0 263.34 ;
   RECT 23.18 263.34 418.0 265.05 ;
   RECT 23.18 265.05 418.0 266.76 ;
   RECT 23.18 266.76 418.0 268.47 ;
   RECT 23.18 268.47 418.0 270.18 ;
   RECT 23.18 270.18 418.0 271.89 ;
   RECT 23.18 271.89 418.0 273.6 ;
   RECT 23.18 273.6 418.0 275.31 ;
   RECT 23.18 275.31 418.0 277.02 ;
   RECT 23.18 277.02 418.0 278.73 ;
   RECT 23.18 278.73 418.0 280.44 ;
   RECT 23.18 280.44 418.0 282.15 ;
   RECT 23.18 282.15 418.0 283.86 ;
   RECT 23.18 283.86 418.0 285.57 ;
   RECT 23.18 285.57 418.0 287.28 ;
   RECT 23.18 287.28 418.0 288.99 ;
   RECT 23.18 288.99 418.0 290.7 ;
   RECT 23.18 290.7 418.0 292.41 ;
   RECT 23.18 292.41 418.0 294.12 ;
   RECT 23.18 294.12 418.0 295.83 ;
  LAYER via3 ;
   RECT 23.18 0.0 418.0 1.71 ;
   RECT 23.18 1.71 418.0 3.42 ;
   RECT 23.18 3.42 418.0 5.13 ;
   RECT 23.18 5.13 418.0 6.84 ;
   RECT 23.18 6.84 418.0 8.55 ;
   RECT 23.18 8.55 418.0 10.26 ;
   RECT 23.18 10.26 418.0 11.97 ;
   RECT 23.18 11.97 418.0 13.68 ;
   RECT 23.18 13.68 418.0 15.39 ;
   RECT 23.18 15.39 418.0 17.1 ;
   RECT 23.18 17.1 418.0 18.81 ;
   RECT 23.18 18.81 418.0 20.52 ;
   RECT 23.18 20.52 418.0 22.23 ;
   RECT 23.18 22.23 418.0 23.94 ;
   RECT 23.18 23.94 418.0 25.65 ;
   RECT 23.18 25.65 418.0 27.36 ;
   RECT 23.18 27.36 418.0 29.07 ;
   RECT 23.18 29.07 418.0 30.78 ;
   RECT 23.18 30.78 418.0 32.49 ;
   RECT 23.18 32.49 418.0 34.2 ;
   RECT 23.18 34.2 418.0 35.91 ;
   RECT 23.18 35.91 418.0 37.62 ;
   RECT 23.18 37.62 418.0 39.33 ;
   RECT 23.18 39.33 418.0 41.04 ;
   RECT 23.18 41.04 418.0 42.75 ;
   RECT 23.18 42.75 418.0 44.46 ;
   RECT 23.18 44.46 418.0 46.17 ;
   RECT 23.18 46.17 418.0 47.88 ;
   RECT 23.18 47.88 418.0 49.59 ;
   RECT 23.18 49.59 418.0 51.3 ;
   RECT 23.18 51.3 418.0 53.01 ;
   RECT 23.18 53.01 418.0 54.72 ;
   RECT 23.18 54.72 418.0 56.43 ;
   RECT 23.18 56.43 418.0 58.14 ;
   RECT 23.18 58.14 418.0 59.85 ;
   RECT 23.18 59.85 418.0 61.56 ;
   RECT 23.18 61.56 418.0 63.27 ;
   RECT 23.18 63.27 418.0 64.98 ;
   RECT 23.18 64.98 418.0 66.69 ;
   RECT 23.18 66.69 418.0 68.4 ;
   RECT 23.18 68.4 418.0 70.11 ;
   RECT 23.18 70.11 418.0 71.82 ;
   RECT 23.18 71.82 418.0 73.53 ;
   RECT 23.18 73.53 418.0 75.24 ;
   RECT 23.18 75.24 418.0 76.95 ;
   RECT 23.18 76.95 418.0 78.66 ;
   RECT 23.18 78.66 418.0 80.37 ;
   RECT 23.18 80.37 418.0 82.08 ;
   RECT 23.18 82.08 418.0 83.79 ;
   RECT 23.18 83.79 418.0 85.5 ;
   RECT 23.18 85.5 418.0 87.21 ;
   RECT 23.18 87.21 418.0 88.92 ;
   RECT 23.18 88.92 418.0 90.63 ;
   RECT 23.18 90.63 418.0 92.34 ;
   RECT 23.18 92.34 418.0 94.05 ;
   RECT 23.18 94.05 418.0 95.76 ;
   RECT 23.18 95.76 418.0 97.47 ;
   RECT 23.18 97.47 418.0 99.18 ;
   RECT 23.18 99.18 418.0 100.89 ;
   RECT 23.18 100.89 418.0 102.6 ;
   RECT 23.18 102.6 418.0 104.31 ;
   RECT 23.18 104.31 418.0 106.02 ;
   RECT 23.18 106.02 418.0 107.73 ;
   RECT 23.18 107.73 418.0 109.44 ;
   RECT 23.18 109.44 418.0 111.15 ;
   RECT 23.18 111.15 418.0 112.86 ;
   RECT 23.18 112.86 418.0 114.57 ;
   RECT 23.18 114.57 418.0 116.28 ;
   RECT 23.18 116.28 418.0 117.99 ;
   RECT 23.18 117.99 418.0 119.7 ;
   RECT 23.18 119.7 418.0 121.41 ;
   RECT 23.18 121.41 418.0 123.12 ;
   RECT 23.18 123.12 418.0 124.83 ;
   RECT 23.18 124.83 418.0 126.54 ;
   RECT 23.18 126.54 418.0 128.25 ;
   RECT 23.18 128.25 418.0 129.96 ;
   RECT 23.18 129.96 418.0 131.67 ;
   RECT 23.18 131.67 418.0 133.38 ;
   RECT 0.0 133.38 418.0 135.09 ;
   RECT 0.0 135.09 418.0 136.8 ;
   RECT 0.0 136.8 418.0 138.51 ;
   RECT 0.0 138.51 418.0 140.22 ;
   RECT 0.0 140.22 418.0 141.93 ;
   RECT 0.0 141.93 418.0 143.64 ;
   RECT 0.0 143.64 418.0 145.35 ;
   RECT 0.0 145.35 418.0 147.06 ;
   RECT 0.0 147.06 418.0 148.77 ;
   RECT 0.0 148.77 418.0 150.48 ;
   RECT 0.0 150.48 418.0 152.19 ;
   RECT 0.0 152.19 418.0 153.9 ;
   RECT 0.0 153.9 418.0 155.61 ;
   RECT 0.0 155.61 418.0 157.32 ;
   RECT 0.0 157.32 418.0 159.03 ;
   RECT 0.0 159.03 418.0 160.74 ;
   RECT 0.0 160.74 418.0 162.45 ;
   RECT 23.18 162.45 418.0 164.16 ;
   RECT 23.18 164.16 418.0 165.87 ;
   RECT 23.18 165.87 418.0 167.58 ;
   RECT 23.18 167.58 418.0 169.29 ;
   RECT 23.18 169.29 418.0 171.0 ;
   RECT 23.18 171.0 418.0 172.71 ;
   RECT 23.18 172.71 418.0 174.42 ;
   RECT 23.18 174.42 418.0 176.13 ;
   RECT 23.18 176.13 418.0 177.84 ;
   RECT 23.18 177.84 418.0 179.55 ;
   RECT 23.18 179.55 418.0 181.26 ;
   RECT 23.18 181.26 418.0 182.97 ;
   RECT 23.18 182.97 418.0 184.68 ;
   RECT 23.18 184.68 418.0 186.39 ;
   RECT 23.18 186.39 418.0 188.1 ;
   RECT 23.18 188.1 418.0 189.81 ;
   RECT 23.18 189.81 418.0 191.52 ;
   RECT 23.18 191.52 418.0 193.23 ;
   RECT 23.18 193.23 418.0 194.94 ;
   RECT 23.18 194.94 418.0 196.65 ;
   RECT 23.18 196.65 418.0 198.36 ;
   RECT 23.18 198.36 418.0 200.07 ;
   RECT 23.18 200.07 418.0 201.78 ;
   RECT 23.18 201.78 418.0 203.49 ;
   RECT 23.18 203.49 418.0 205.2 ;
   RECT 23.18 205.2 418.0 206.91 ;
   RECT 23.18 206.91 418.0 208.62 ;
   RECT 23.18 208.62 418.0 210.33 ;
   RECT 23.18 210.33 418.0 212.04 ;
   RECT 23.18 212.04 418.0 213.75 ;
   RECT 23.18 213.75 418.0 215.46 ;
   RECT 23.18 215.46 418.0 217.17 ;
   RECT 23.18 217.17 418.0 218.88 ;
   RECT 23.18 218.88 418.0 220.59 ;
   RECT 23.18 220.59 418.0 222.3 ;
   RECT 23.18 222.3 418.0 224.01 ;
   RECT 23.18 224.01 418.0 225.72 ;
   RECT 23.18 225.72 418.0 227.43 ;
   RECT 23.18 227.43 418.0 229.14 ;
   RECT 23.18 229.14 418.0 230.85 ;
   RECT 23.18 230.85 418.0 232.56 ;
   RECT 23.18 232.56 418.0 234.27 ;
   RECT 23.18 234.27 418.0 235.98 ;
   RECT 23.18 235.98 418.0 237.69 ;
   RECT 23.18 237.69 418.0 239.4 ;
   RECT 23.18 239.4 418.0 241.11 ;
   RECT 23.18 241.11 418.0 242.82 ;
   RECT 23.18 242.82 418.0 244.53 ;
   RECT 23.18 244.53 418.0 246.24 ;
   RECT 23.18 246.24 418.0 247.95 ;
   RECT 23.18 247.95 418.0 249.66 ;
   RECT 23.18 249.66 418.0 251.37 ;
   RECT 23.18 251.37 418.0 253.08 ;
   RECT 23.18 253.08 418.0 254.79 ;
   RECT 23.18 254.79 418.0 256.5 ;
   RECT 23.18 256.5 418.0 258.21 ;
   RECT 23.18 258.21 418.0 259.92 ;
   RECT 23.18 259.92 418.0 261.63 ;
   RECT 23.18 261.63 418.0 263.34 ;
   RECT 23.18 263.34 418.0 265.05 ;
   RECT 23.18 265.05 418.0 266.76 ;
   RECT 23.18 266.76 418.0 268.47 ;
   RECT 23.18 268.47 418.0 270.18 ;
   RECT 23.18 270.18 418.0 271.89 ;
   RECT 23.18 271.89 418.0 273.6 ;
   RECT 23.18 273.6 418.0 275.31 ;
   RECT 23.18 275.31 418.0 277.02 ;
   RECT 23.18 277.02 418.0 278.73 ;
   RECT 23.18 278.73 418.0 280.44 ;
   RECT 23.18 280.44 418.0 282.15 ;
   RECT 23.18 282.15 418.0 283.86 ;
   RECT 23.18 283.86 418.0 285.57 ;
   RECT 23.18 285.57 418.0 287.28 ;
   RECT 23.18 287.28 418.0 288.99 ;
   RECT 23.18 288.99 418.0 290.7 ;
   RECT 23.18 290.7 418.0 292.41 ;
   RECT 23.18 292.41 418.0 294.12 ;
   RECT 23.18 294.12 418.0 295.83 ;
  LAYER metal4 ;
   RECT 23.18 0.0 418.0 1.71 ;
   RECT 23.18 1.71 418.0 3.42 ;
   RECT 23.18 3.42 418.0 5.13 ;
   RECT 23.18 5.13 418.0 6.84 ;
   RECT 23.18 6.84 418.0 8.55 ;
   RECT 23.18 8.55 418.0 10.26 ;
   RECT 23.18 10.26 418.0 11.97 ;
   RECT 23.18 11.97 418.0 13.68 ;
   RECT 23.18 13.68 418.0 15.39 ;
   RECT 23.18 15.39 418.0 17.1 ;
   RECT 23.18 17.1 418.0 18.81 ;
   RECT 23.18 18.81 418.0 20.52 ;
   RECT 23.18 20.52 418.0 22.23 ;
   RECT 23.18 22.23 418.0 23.94 ;
   RECT 23.18 23.94 418.0 25.65 ;
   RECT 23.18 25.65 418.0 27.36 ;
   RECT 23.18 27.36 418.0 29.07 ;
   RECT 23.18 29.07 418.0 30.78 ;
   RECT 23.18 30.78 418.0 32.49 ;
   RECT 23.18 32.49 418.0 34.2 ;
   RECT 23.18 34.2 418.0 35.91 ;
   RECT 23.18 35.91 418.0 37.62 ;
   RECT 23.18 37.62 418.0 39.33 ;
   RECT 23.18 39.33 418.0 41.04 ;
   RECT 23.18 41.04 418.0 42.75 ;
   RECT 23.18 42.75 418.0 44.46 ;
   RECT 23.18 44.46 418.0 46.17 ;
   RECT 23.18 46.17 418.0 47.88 ;
   RECT 23.18 47.88 418.0 49.59 ;
   RECT 23.18 49.59 418.0 51.3 ;
   RECT 23.18 51.3 418.0 53.01 ;
   RECT 23.18 53.01 418.0 54.72 ;
   RECT 23.18 54.72 418.0 56.43 ;
   RECT 23.18 56.43 418.0 58.14 ;
   RECT 23.18 58.14 418.0 59.85 ;
   RECT 23.18 59.85 418.0 61.56 ;
   RECT 23.18 61.56 418.0 63.27 ;
   RECT 23.18 63.27 418.0 64.98 ;
   RECT 23.18 64.98 418.0 66.69 ;
   RECT 23.18 66.69 418.0 68.4 ;
   RECT 23.18 68.4 418.0 70.11 ;
   RECT 23.18 70.11 418.0 71.82 ;
   RECT 23.18 71.82 418.0 73.53 ;
   RECT 23.18 73.53 418.0 75.24 ;
   RECT 23.18 75.24 418.0 76.95 ;
   RECT 23.18 76.95 418.0 78.66 ;
   RECT 23.18 78.66 418.0 80.37 ;
   RECT 23.18 80.37 418.0 82.08 ;
   RECT 23.18 82.08 418.0 83.79 ;
   RECT 23.18 83.79 418.0 85.5 ;
   RECT 23.18 85.5 418.0 87.21 ;
   RECT 23.18 87.21 418.0 88.92 ;
   RECT 23.18 88.92 418.0 90.63 ;
   RECT 23.18 90.63 418.0 92.34 ;
   RECT 23.18 92.34 418.0 94.05 ;
   RECT 23.18 94.05 418.0 95.76 ;
   RECT 23.18 95.76 418.0 97.47 ;
   RECT 23.18 97.47 418.0 99.18 ;
   RECT 23.18 99.18 418.0 100.89 ;
   RECT 23.18 100.89 418.0 102.6 ;
   RECT 23.18 102.6 418.0 104.31 ;
   RECT 23.18 104.31 418.0 106.02 ;
   RECT 23.18 106.02 418.0 107.73 ;
   RECT 23.18 107.73 418.0 109.44 ;
   RECT 23.18 109.44 418.0 111.15 ;
   RECT 23.18 111.15 418.0 112.86 ;
   RECT 23.18 112.86 418.0 114.57 ;
   RECT 23.18 114.57 418.0 116.28 ;
   RECT 23.18 116.28 418.0 117.99 ;
   RECT 23.18 117.99 418.0 119.7 ;
   RECT 23.18 119.7 418.0 121.41 ;
   RECT 23.18 121.41 418.0 123.12 ;
   RECT 23.18 123.12 418.0 124.83 ;
   RECT 23.18 124.83 418.0 126.54 ;
   RECT 23.18 126.54 418.0 128.25 ;
   RECT 23.18 128.25 418.0 129.96 ;
   RECT 23.18 129.96 418.0 131.67 ;
   RECT 23.18 131.67 418.0 133.38 ;
   RECT 0.0 133.38 418.0 135.09 ;
   RECT 0.0 135.09 418.0 136.8 ;
   RECT 0.0 136.8 418.0 138.51 ;
   RECT 0.0 138.51 418.0 140.22 ;
   RECT 0.0 140.22 418.0 141.93 ;
   RECT 0.0 141.93 418.0 143.64 ;
   RECT 0.0 143.64 418.0 145.35 ;
   RECT 0.0 145.35 418.0 147.06 ;
   RECT 0.0 147.06 418.0 148.77 ;
   RECT 0.0 148.77 418.0 150.48 ;
   RECT 0.0 150.48 418.0 152.19 ;
   RECT 0.0 152.19 418.0 153.9 ;
   RECT 0.0 153.9 418.0 155.61 ;
   RECT 0.0 155.61 418.0 157.32 ;
   RECT 0.0 157.32 418.0 159.03 ;
   RECT 0.0 159.03 418.0 160.74 ;
   RECT 0.0 160.74 418.0 162.45 ;
   RECT 23.18 162.45 418.0 164.16 ;
   RECT 23.18 164.16 418.0 165.87 ;
   RECT 23.18 165.87 418.0 167.58 ;
   RECT 23.18 167.58 418.0 169.29 ;
   RECT 23.18 169.29 418.0 171.0 ;
   RECT 23.18 171.0 418.0 172.71 ;
   RECT 23.18 172.71 418.0 174.42 ;
   RECT 23.18 174.42 418.0 176.13 ;
   RECT 23.18 176.13 418.0 177.84 ;
   RECT 23.18 177.84 418.0 179.55 ;
   RECT 23.18 179.55 418.0 181.26 ;
   RECT 23.18 181.26 418.0 182.97 ;
   RECT 23.18 182.97 418.0 184.68 ;
   RECT 23.18 184.68 418.0 186.39 ;
   RECT 23.18 186.39 418.0 188.1 ;
   RECT 23.18 188.1 418.0 189.81 ;
   RECT 23.18 189.81 418.0 191.52 ;
   RECT 23.18 191.52 418.0 193.23 ;
   RECT 23.18 193.23 418.0 194.94 ;
   RECT 23.18 194.94 418.0 196.65 ;
   RECT 23.18 196.65 418.0 198.36 ;
   RECT 23.18 198.36 418.0 200.07 ;
   RECT 23.18 200.07 418.0 201.78 ;
   RECT 23.18 201.78 418.0 203.49 ;
   RECT 23.18 203.49 418.0 205.2 ;
   RECT 23.18 205.2 418.0 206.91 ;
   RECT 23.18 206.91 418.0 208.62 ;
   RECT 23.18 208.62 418.0 210.33 ;
   RECT 23.18 210.33 418.0 212.04 ;
   RECT 23.18 212.04 418.0 213.75 ;
   RECT 23.18 213.75 418.0 215.46 ;
   RECT 23.18 215.46 418.0 217.17 ;
   RECT 23.18 217.17 418.0 218.88 ;
   RECT 23.18 218.88 418.0 220.59 ;
   RECT 23.18 220.59 418.0 222.3 ;
   RECT 23.18 222.3 418.0 224.01 ;
   RECT 23.18 224.01 418.0 225.72 ;
   RECT 23.18 225.72 418.0 227.43 ;
   RECT 23.18 227.43 418.0 229.14 ;
   RECT 23.18 229.14 418.0 230.85 ;
   RECT 23.18 230.85 418.0 232.56 ;
   RECT 23.18 232.56 418.0 234.27 ;
   RECT 23.18 234.27 418.0 235.98 ;
   RECT 23.18 235.98 418.0 237.69 ;
   RECT 23.18 237.69 418.0 239.4 ;
   RECT 23.18 239.4 418.0 241.11 ;
   RECT 23.18 241.11 418.0 242.82 ;
   RECT 23.18 242.82 418.0 244.53 ;
   RECT 23.18 244.53 418.0 246.24 ;
   RECT 23.18 246.24 418.0 247.95 ;
   RECT 23.18 247.95 418.0 249.66 ;
   RECT 23.18 249.66 418.0 251.37 ;
   RECT 23.18 251.37 418.0 253.08 ;
   RECT 23.18 253.08 418.0 254.79 ;
   RECT 23.18 254.79 418.0 256.5 ;
   RECT 23.18 256.5 418.0 258.21 ;
   RECT 23.18 258.21 418.0 259.92 ;
   RECT 23.18 259.92 418.0 261.63 ;
   RECT 23.18 261.63 418.0 263.34 ;
   RECT 23.18 263.34 418.0 265.05 ;
   RECT 23.18 265.05 418.0 266.76 ;
   RECT 23.18 266.76 418.0 268.47 ;
   RECT 23.18 268.47 418.0 270.18 ;
   RECT 23.18 270.18 418.0 271.89 ;
   RECT 23.18 271.89 418.0 273.6 ;
   RECT 23.18 273.6 418.0 275.31 ;
   RECT 23.18 275.31 418.0 277.02 ;
   RECT 23.18 277.02 418.0 278.73 ;
   RECT 23.18 278.73 418.0 280.44 ;
   RECT 23.18 280.44 418.0 282.15 ;
   RECT 23.18 282.15 418.0 283.86 ;
   RECT 23.18 283.86 418.0 285.57 ;
   RECT 23.18 285.57 418.0 287.28 ;
   RECT 23.18 287.28 418.0 288.99 ;
   RECT 23.18 288.99 418.0 290.7 ;
   RECT 23.18 290.7 418.0 292.41 ;
   RECT 23.18 292.41 418.0 294.12 ;
   RECT 23.18 294.12 418.0 295.83 ;
 END
END block_1100x1557_168

MACRO block_341x369_78
 CLASS BLOCK ;
 FOREIGN block_341x369_78 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 129.58 BY 70.11 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 20.235 126.445 20.805 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 26.695 126.445 27.265 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 6.935 3.325 7.505 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 7.695 3.325 8.265 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 9.215 3.325 9.785 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 10.735 3.325 11.305 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 11.495 3.325 12.065 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 13.015 3.325 13.585 ;
  END
 END o7
 PIN o8
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 13.395 4.085 13.965 ;
  END
 END o8
 PIN o9
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 13.775 3.325 14.345 ;
  END
 END o9
 PIN o10
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 15.295 3.325 15.865 ;
  END
 END o10
 PIN o11
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 16.055 3.325 16.625 ;
  END
 END o11
 PIN o12
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 12.635 4.085 13.205 ;
  END
 END o12
 PIN o13
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 19.855 3.325 20.425 ;
  END
 END o13
 PIN o14
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 20.615 3.325 21.185 ;
  END
 END o14
 PIN o15
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 21.375 3.325 21.945 ;
  END
 END o15
 PIN o16
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 22.135 3.325 22.705 ;
  END
 END o16
 PIN o17
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 18.335 3.325 18.905 ;
  END
 END o17
 PIN o18
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 25.935 3.325 26.505 ;
  END
 END o18
 PIN o19
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 26.695 3.325 27.265 ;
  END
 END o19
 PIN o20
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 27.455 3.325 28.025 ;
  END
 END o20
 PIN o21
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 28.975 3.325 29.545 ;
  END
 END o21
 PIN o22
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 25.175 3.325 25.745 ;
  END
 END o22
 PIN o23
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 32.015 3.325 32.585 ;
  END
 END o23
 PIN o24
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 33.535 3.325 34.105 ;
  END
 END o24
 PIN o25
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 34.295 3.325 34.865 ;
  END
 END o25
 PIN o26
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 35.055 3.325 35.625 ;
  END
 END o26
 PIN o27
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 31.255 3.325 31.825 ;
  END
 END o27
 PIN o28
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 38.095 126.445 38.665 ;
  END
 END o28
 PIN o29
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 38.855 126.445 39.425 ;
  END
 END o29
 PIN o30
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 39.615 126.445 40.185 ;
  END
 END o30
 PIN o31
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 42.655 126.445 43.225 ;
  END
 END o31
 PIN o32
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 29.735 126.445 30.305 ;
  END
 END o32
 PIN o33
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 21.755 126.445 22.325 ;
  END
 END o33
 PIN o34
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 31.255 126.445 31.825 ;
  END
 END o34
 PIN o35
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 32.015 126.445 32.585 ;
  END
 END o35
 PIN o36
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 33.535 126.445 34.105 ;
  END
 END o36
 PIN o37
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 34.295 126.445 34.865 ;
  END
 END o37
 PIN o38
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 35.055 126.445 35.625 ;
  END
 END o38
 PIN o39
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 30.495 126.445 31.065 ;
  END
 END o39
 PIN o40
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 28.975 126.445 29.545 ;
  END
 END o40
 PIN o41
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 41.135 3.325 41.705 ;
  END
 END o41
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 35.815 126.445 36.385 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 43.035 125.685 43.605 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 32.395 125.685 32.965 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 35.435 125.685 36.005 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 36.955 126.445 37.525 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 36.575 125.685 37.145 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 33.915 125.685 34.485 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 30.115 125.685 30.685 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 8.455 3.325 9.025 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 25.935 126.445 26.505 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 25.175 126.445 25.745 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 24.415 126.445 24.985 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 34.675 125.685 35.245 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 30.875 125.685 31.445 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 40.755 126.445 41.325 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 40.375 3.325 40.945 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 27.455 126.445 28.025 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 38.475 125.685 39.045 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 39.995 125.685 40.565 ;
  END
 END i18
 PIN i19
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 39.235 125.685 39.805 ;
  END
 END i19
 PIN i20
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 124.355 40.375 124.925 40.945 ;
  END
 END i20
 PIN i21
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 8.455 126.445 9.025 ;
  END
 END i21
 PIN i22
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 9.215 126.445 9.785 ;
  END
 END i22
 PIN i23
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 10.735 126.445 11.305 ;
  END
 END i23
 PIN i24
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 11.495 126.445 12.065 ;
  END
 END i24
 PIN i25
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 12.255 126.445 12.825 ;
  END
 END i25
 PIN i26
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 13.015 126.445 13.585 ;
  END
 END i26
 PIN i27
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 8.075 125.685 8.645 ;
  END
 END i27
 PIN i28
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 7.695 126.445 8.265 ;
  END
 END i28
 PIN i29
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 7.315 125.685 7.885 ;
  END
 END i29
 PIN i30
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 6.935 126.445 7.505 ;
  END
 END i30
 PIN i31
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.115 6.555 125.685 7.125 ;
  END
 END i31
 PIN i32
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 13.775 126.445 14.345 ;
  END
 END i32
 PIN i33
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 15.295 126.445 15.865 ;
  END
 END i33
 PIN i34
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 16.055 126.445 16.625 ;
  END
 END i34
 PIN i35
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 125.875 16.815 126.445 17.385 ;
  END
 END i35
 OBS
  LAYER metal1 ;
   RECT 0 0 129.58 70.11 ;
  LAYER via1 ;
   RECT 0 0 129.58 70.11 ;
  LAYER metal2 ;
   RECT 0 0 129.58 70.11 ;
  LAYER via2 ;
   RECT 0 0 129.58 70.11 ;
  LAYER metal3 ;
   RECT 0 0 129.58 70.11 ;
  LAYER via3 ;
   RECT 0 0 129.58 70.11 ;
  LAYER metal4 ;
   RECT 0 0 129.58 70.11 ;
 END
END block_341x369_78

MACRO block_315x981_72
 CLASS BLOCK ;
 FOREIGN block_315x981_72 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 119.7 BY 186.39 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 131.765 9.785 132.335 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 137.465 9.785 138.035 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 143.355 9.785 143.925 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 149.055 9.785 149.625 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 154.755 9.785 155.325 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 160.455 9.785 161.025 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 166.345 9.785 166.915 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 172.045 9.785 172.615 ;
  END
 END o7
 PIN o8
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 8.265 9.785 8.835 ;
  END
 END o8
 PIN o9
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 13.965 9.785 14.535 ;
  END
 END o9
 PIN o10
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 19.855 9.785 20.425 ;
  END
 END o10
 PIN o11
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 25.555 9.785 26.125 ;
  END
 END o11
 PIN o12
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 31.255 9.785 31.825 ;
  END
 END o12
 PIN o13
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 36.955 9.785 37.525 ;
  END
 END o13
 PIN o14
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 42.845 9.785 43.415 ;
  END
 END o14
 PIN o15
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 177.745 9.785 178.315 ;
  END
 END o15
 PIN o16
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 48.545 9.785 49.115 ;
  END
 END o16
 PIN o17
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 54.245 9.785 54.815 ;
  END
 END o17
 PIN o18
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 59.945 9.785 60.515 ;
  END
 END o18
 PIN o19
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 65.835 9.785 66.405 ;
  END
 END o19
 PIN o20
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 71.535 9.785 72.105 ;
  END
 END o20
 PIN o21
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 77.235 9.785 77.805 ;
  END
 END o21
 PIN o22
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 108.775 9.785 109.345 ;
  END
 END o22
 PIN o23
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 114.475 9.785 115.045 ;
  END
 END o23
 PIN o24
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 120.365 9.785 120.935 ;
  END
 END o24
 PIN o25
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 126.065 9.785 126.635 ;
  END
 END o25
 PIN o26
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 183.445 9.785 184.015 ;
  END
 END o26
 PIN o27
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 2.565 9.785 3.135 ;
  END
 END o27
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 94.525 118.465 95.095 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 85.025 118.465 85.595 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 111.815 85.215 112.385 85.785 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 86.355 118.465 86.925 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 87.685 118.465 88.255 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.135 88.255 117.705 88.825 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 85.975 9.785 86.545 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 101.745 118.465 102.315 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 91.865 118.465 92.435 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 93.005 118.465 93.575 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 93.005 9.785 93.575 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 8.455 99.655 9.025 100.225 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 96.615 9.785 97.185 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.135 94.905 117.705 95.475 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 96.805 118.465 97.375 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.135 97.185 117.705 97.755 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 183.065 118.465 183.635 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 125.685 118.465 126.255 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 119.795 118.465 120.365 ;
  END
 END i18
 PIN i19
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 114.095 118.465 114.665 ;
  END
 END i19
 PIN i20
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 108.395 118.465 108.965 ;
  END
 END i20
 PIN i21
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 77.615 118.465 78.185 ;
  END
 END i21
 PIN i22
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 71.915 118.465 72.485 ;
  END
 END i22
 PIN i23
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 66.215 118.465 66.785 ;
  END
 END i23
 PIN i24
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 60.515 118.465 61.085 ;
  END
 END i24
 PIN i25
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 54.625 118.465 55.195 ;
  END
 END i25
 PIN i26
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 48.925 118.465 49.495 ;
  END
 END i26
 PIN i27
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 177.365 118.465 177.935 ;
  END
 END i27
 PIN i28
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 43.225 118.465 43.795 ;
  END
 END i28
 PIN i29
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 37.525 118.465 38.095 ;
  END
 END i29
 PIN i30
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 31.635 118.465 32.205 ;
  END
 END i30
 PIN i31
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 25.935 118.465 26.505 ;
  END
 END i31
 PIN i32
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 20.235 118.465 20.805 ;
  END
 END i32
 PIN i33
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 14.535 118.465 15.105 ;
  END
 END i33
 PIN i34
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 8.645 118.465 9.215 ;
  END
 END i34
 PIN i35
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 2.945 118.465 3.515 ;
  END
 END i35
 PIN i36
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 171.665 118.465 172.235 ;
  END
 END i36
 PIN i37
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 165.775 118.465 166.345 ;
  END
 END i37
 PIN i38
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 160.075 118.465 160.645 ;
  END
 END i38
 PIN i39
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 154.375 118.465 154.945 ;
  END
 END i39
 PIN i40
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 148.675 118.465 149.245 ;
  END
 END i40
 PIN i41
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 142.785 118.465 143.355 ;
  END
 END i41
 PIN i42
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 137.085 118.465 137.655 ;
  END
 END i42
 PIN i43
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 131.385 118.465 131.955 ;
  END
 END i43
 OBS
  LAYER metal1 ;
   RECT 0 0 119.7 186.39 ;
  LAYER via1 ;
   RECT 0 0 119.7 186.39 ;
  LAYER metal2 ;
   RECT 0 0 119.7 186.39 ;
  LAYER via2 ;
   RECT 0 0 119.7 186.39 ;
  LAYER metal3 ;
   RECT 0 0 119.7 186.39 ;
  LAYER via3 ;
   RECT 0 0 119.7 186.39 ;
  LAYER metal4 ;
   RECT 0 0 119.7 186.39 ;
 END
END block_315x981_72

MACRO block_535x756_102
 CLASS BLOCK ;
 FOREIGN block_535x756_102 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 203.3 BY 143.64 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 107.445 56.525 108.015 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 97.945 56.525 98.515 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 88.445 56.525 89.015 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 78.945 56.525 79.515 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 69.445 56.525 70.015 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 50.445 56.525 51.015 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 59.945 56.525 60.515 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 40.945 56.525 41.515 ;
  END
 END o7
 PIN o8
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 25.555 3.705 26.125 ;
  END
 END o8
 PIN o9
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 116.945 56.525 117.515 ;
  END
 END o9
 PIN o10
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 37.715 56.525 38.285 ;
  END
 END o10
 PIN o11
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 47.215 56.525 47.785 ;
  END
 END o11
 PIN o12
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 56.715 56.525 57.285 ;
  END
 END o12
 PIN o13
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 66.215 56.525 66.785 ;
  END
 END o13
 PIN o14
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 75.715 56.525 76.285 ;
  END
 END o14
 PIN o15
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 85.215 56.525 85.785 ;
  END
 END o15
 PIN o16
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 94.715 56.525 95.285 ;
  END
 END o16
 PIN o17
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 104.215 56.525 104.785 ;
  END
 END o17
 PIN o18
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 113.715 56.525 114.285 ;
  END
 END o18
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 18.145 3.705 18.715 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 16.435 3.705 17.005 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 19.095 3.705 19.665 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 13.395 3.705 13.965 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 16.055 4.465 16.625 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 23.275 3.705 23.845 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 4.655 3.705 5.225 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 5.605 3.705 6.175 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 6.555 3.705 7.125 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 82.555 56.525 83.125 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 101.555 56.525 102.125 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 92.055 56.525 92.625 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 73.055 56.525 73.625 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 63.555 56.525 64.125 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 54.055 56.525 54.625 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 44.555 56.525 45.125 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 35.055 56.525 35.625 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 111.055 56.525 111.625 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 0.855 3.705 1.425 ;
  END
 END i18
 PIN i19
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 26.125 4.465 26.695 ;
  END
 END i19
 PIN i20
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 118.465 56.525 119.035 ;
  END
 END i20
 PIN i21
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 56.715 118.845 57.285 119.415 ;
  END
 END i21
 PIN i22
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 120.555 56.525 121.125 ;
  END
 END i22
 PIN i23
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 119.225 56.525 119.795 ;
  END
 END i23
 PIN i24
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 56.715 119.795 57.285 120.365 ;
  END
 END i24
 PIN i25
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 30.495 3.705 31.065 ;
  END
 END i25
 PIN i26
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 28.975 3.705 29.545 ;
  END
 END i26
 PIN i27
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 2.375 3.705 2.945 ;
  END
 END i27
 PIN i28
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 1.805 4.465 2.375 ;
  END
 END i28
 PIN i29
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 29.925 4.465 30.495 ;
  END
 END i29
 PIN i30
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 28.025 3.705 28.595 ;
  END
 END i30
 PIN i31
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 2.755 4.465 3.325 ;
  END
 END i31
 PIN i32
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 4.275 4.465 4.845 ;
  END
 END i32
 PIN i33
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 3.705 3.705 4.275 ;
  END
 END i33
 PIN i34
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 4.655 29.545 5.225 30.115 ;
  END
 END i34
 PIN i35
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 13.775 4.465 14.345 ;
  END
 END i35
 PIN i36
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 18.525 4.465 19.095 ;
  END
 END i36
 PIN i37
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 17.575 4.465 18.145 ;
  END
 END i37
 PIN i38
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 23.655 4.465 24.225 ;
  END
 END i38
 PIN i39
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 24.225 3.705 24.795 ;
  END
 END i39
 PIN i40
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 5.225 4.465 5.795 ;
  END
 END i40
 PIN i41
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 6.175 4.465 6.745 ;
  END
 END i41
 PIN i42
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 7.125 4.465 7.695 ;
  END
 END i42
 PIN i43
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 10.925 3.705 11.495 ;
  END
 END i43
 PIN i44
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 26.505 3.705 27.075 ;
  END
 END i44
 PIN i45
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 4.655 1.425 5.225 1.995 ;
  END
 END i45
 PIN i46
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 33.725 56.525 34.295 ;
  END
 END i46
 PIN i47
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 43.225 56.525 43.795 ;
  END
 END i47
 PIN i48
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 52.725 56.525 53.295 ;
  END
 END i48
 PIN i49
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 62.225 56.525 62.795 ;
  END
 END i49
 PIN i50
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 71.725 56.525 72.295 ;
  END
 END i50
 PIN i51
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 81.225 56.525 81.795 ;
  END
 END i51
 PIN i52
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 90.725 56.525 91.295 ;
  END
 END i52
 PIN i53
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 100.225 56.525 100.795 ;
  END
 END i53
 PIN i54
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 109.725 56.525 110.295 ;
  END
 END i54
 PIN i55
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 38.855 56.525 39.425 ;
  END
 END i55
 PIN i56
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 48.355 56.525 48.925 ;
  END
 END i56
 PIN i57
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 57.855 56.525 58.425 ;
  END
 END i57
 PIN i58
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 67.355 56.525 67.925 ;
  END
 END i58
 PIN i59
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 76.855 56.525 77.425 ;
  END
 END i59
 PIN i60
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 86.355 56.525 86.925 ;
  END
 END i60
 PIN i61
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 95.855 56.525 96.425 ;
  END
 END i61
 PIN i62
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 105.355 56.525 105.925 ;
  END
 END i62
 PIN i63
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 114.855 56.525 115.425 ;
  END
 END i63
 PIN i64
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 56.715 120.935 57.285 121.505 ;
  END
 END i64
 PIN i65
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 39.805 56.525 40.375 ;
  END
 END i65
 PIN i66
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 49.305 56.525 49.875 ;
  END
 END i66
 PIN i67
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 58.805 56.525 59.375 ;
  END
 END i67
 PIN i68
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 68.305 56.525 68.875 ;
  END
 END i68
 PIN i69
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 77.805 56.525 78.375 ;
  END
 END i69
 PIN i70
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 87.305 56.525 87.875 ;
  END
 END i70
 PIN i71
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 96.805 56.525 97.375 ;
  END
 END i71
 PIN i72
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 106.305 56.525 106.875 ;
  END
 END i72
 PIN i73
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 55.955 115.805 56.525 116.375 ;
  END
 END i73
 PIN i74
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 56.715 34.105 57.285 34.675 ;
  END
 END i74
 PIN i75
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 56.715 43.605 57.285 44.175 ;
  END
 END i75
 PIN i76
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 56.715 53.105 57.285 53.675 ;
  END
 END i76
 PIN i77
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 56.715 62.605 57.285 63.175 ;
  END
 END i77
 PIN i78
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 56.715 72.105 57.285 72.675 ;
  END
 END i78
 PIN i79
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 56.715 81.605 57.285 82.175 ;
  END
 END i79
 PIN i80
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 56.715 91.105 57.285 91.675 ;
  END
 END i80
 PIN i81
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 56.715 100.605 57.285 101.175 ;
  END
 END i81
 PIN i82
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 56.715 110.105 57.285 110.675 ;
  END
 END i82
 OBS
  LAYER metal1 ;
   RECT 0.0 0.0 203.3 1.71 ;
   RECT 0.0 1.71 203.3 3.42 ;
   RECT 0.0 3.42 203.3 5.13 ;
   RECT 0.0 5.13 203.3 6.84 ;
   RECT 0.0 6.84 203.3 8.55 ;
   RECT 0.0 8.55 203.3 10.26 ;
   RECT 0.0 10.26 203.3 11.97 ;
   RECT 0.0 11.97 203.3 13.68 ;
   RECT 0.0 13.68 203.3 15.39 ;
   RECT 0.0 15.39 203.3 17.1 ;
   RECT 0.0 17.1 203.3 18.81 ;
   RECT 0.0 18.81 203.3 20.52 ;
   RECT 0.0 20.52 203.3 22.23 ;
   RECT 0.0 22.23 203.3 23.94 ;
   RECT 0.0 23.94 203.3 25.65 ;
   RECT 0.0 25.65 203.3 27.36 ;
   RECT 0.0 27.36 203.3 29.07 ;
   RECT 0.0 29.07 203.3 30.78 ;
   RECT 0.0 30.78 203.3 32.49 ;
   RECT 0.0 32.49 203.3 34.2 ;
   RECT 52.82 34.2 203.3 35.91 ;
   RECT 52.82 35.91 203.3 37.62 ;
   RECT 52.82 37.62 203.3 39.33 ;
   RECT 52.82 39.33 203.3 41.04 ;
   RECT 52.82 41.04 203.3 42.75 ;
   RECT 52.82 42.75 203.3 44.46 ;
   RECT 52.82 44.46 203.3 46.17 ;
   RECT 52.82 46.17 203.3 47.88 ;
   RECT 52.82 47.88 203.3 49.59 ;
   RECT 52.82 49.59 203.3 51.3 ;
   RECT 52.82 51.3 203.3 53.01 ;
   RECT 52.82 53.01 203.3 54.72 ;
   RECT 52.82 54.72 203.3 56.43 ;
   RECT 52.82 56.43 203.3 58.14 ;
   RECT 52.82 58.14 203.3 59.85 ;
   RECT 52.82 59.85 203.3 61.56 ;
   RECT 52.82 61.56 203.3 63.27 ;
   RECT 52.82 63.27 203.3 64.98 ;
   RECT 52.82 64.98 203.3 66.69 ;
   RECT 52.82 66.69 203.3 68.4 ;
   RECT 52.82 68.4 203.3 70.11 ;
   RECT 52.82 70.11 203.3 71.82 ;
   RECT 52.82 71.82 203.3 73.53 ;
   RECT 52.82 73.53 203.3 75.24 ;
   RECT 52.82 75.24 203.3 76.95 ;
   RECT 52.82 76.95 203.3 78.66 ;
   RECT 52.82 78.66 203.3 80.37 ;
   RECT 52.82 80.37 203.3 82.08 ;
   RECT 52.82 82.08 203.3 83.79 ;
   RECT 52.82 83.79 203.3 85.5 ;
   RECT 52.82 85.5 203.3 87.21 ;
   RECT 52.82 87.21 203.3 88.92 ;
   RECT 52.82 88.92 203.3 90.63 ;
   RECT 52.82 90.63 203.3 92.34 ;
   RECT 52.82 92.34 203.3 94.05 ;
   RECT 52.82 94.05 203.3 95.76 ;
   RECT 52.82 95.76 203.3 97.47 ;
   RECT 52.82 97.47 203.3 99.18 ;
   RECT 52.82 99.18 203.3 100.89 ;
   RECT 52.82 100.89 203.3 102.6 ;
   RECT 52.82 102.6 203.3 104.31 ;
   RECT 52.82 104.31 203.3 106.02 ;
   RECT 52.82 106.02 203.3 107.73 ;
   RECT 52.82 107.73 203.3 109.44 ;
   RECT 52.82 109.44 203.3 111.15 ;
   RECT 52.82 111.15 203.3 112.86 ;
   RECT 52.82 112.86 203.3 114.57 ;
   RECT 52.82 114.57 203.3 116.28 ;
   RECT 52.82 116.28 203.3 117.99 ;
   RECT 52.82 117.99 203.3 119.7 ;
   RECT 52.82 119.7 203.3 121.41 ;
   RECT 52.82 121.41 203.3 123.12 ;
   RECT 52.82 123.12 203.3 124.83 ;
   RECT 52.82 124.83 203.3 126.54 ;
   RECT 52.82 126.54 203.3 128.25 ;
   RECT 52.82 128.25 203.3 129.96 ;
   RECT 52.82 129.96 203.3 131.67 ;
   RECT 52.82 131.67 203.3 133.38 ;
   RECT 52.82 133.38 203.3 135.09 ;
   RECT 52.82 135.09 203.3 136.8 ;
   RECT 52.82 136.8 203.3 138.51 ;
   RECT 52.82 138.51 203.3 140.22 ;
   RECT 52.82 140.22 203.3 141.93 ;
   RECT 52.82 141.93 203.3 143.64 ;
  LAYER via1 ;
   RECT 0.0 0.0 203.3 1.71 ;
   RECT 0.0 1.71 203.3 3.42 ;
   RECT 0.0 3.42 203.3 5.13 ;
   RECT 0.0 5.13 203.3 6.84 ;
   RECT 0.0 6.84 203.3 8.55 ;
   RECT 0.0 8.55 203.3 10.26 ;
   RECT 0.0 10.26 203.3 11.97 ;
   RECT 0.0 11.97 203.3 13.68 ;
   RECT 0.0 13.68 203.3 15.39 ;
   RECT 0.0 15.39 203.3 17.1 ;
   RECT 0.0 17.1 203.3 18.81 ;
   RECT 0.0 18.81 203.3 20.52 ;
   RECT 0.0 20.52 203.3 22.23 ;
   RECT 0.0 22.23 203.3 23.94 ;
   RECT 0.0 23.94 203.3 25.65 ;
   RECT 0.0 25.65 203.3 27.36 ;
   RECT 0.0 27.36 203.3 29.07 ;
   RECT 0.0 29.07 203.3 30.78 ;
   RECT 0.0 30.78 203.3 32.49 ;
   RECT 0.0 32.49 203.3 34.2 ;
   RECT 52.82 34.2 203.3 35.91 ;
   RECT 52.82 35.91 203.3 37.62 ;
   RECT 52.82 37.62 203.3 39.33 ;
   RECT 52.82 39.33 203.3 41.04 ;
   RECT 52.82 41.04 203.3 42.75 ;
   RECT 52.82 42.75 203.3 44.46 ;
   RECT 52.82 44.46 203.3 46.17 ;
   RECT 52.82 46.17 203.3 47.88 ;
   RECT 52.82 47.88 203.3 49.59 ;
   RECT 52.82 49.59 203.3 51.3 ;
   RECT 52.82 51.3 203.3 53.01 ;
   RECT 52.82 53.01 203.3 54.72 ;
   RECT 52.82 54.72 203.3 56.43 ;
   RECT 52.82 56.43 203.3 58.14 ;
   RECT 52.82 58.14 203.3 59.85 ;
   RECT 52.82 59.85 203.3 61.56 ;
   RECT 52.82 61.56 203.3 63.27 ;
   RECT 52.82 63.27 203.3 64.98 ;
   RECT 52.82 64.98 203.3 66.69 ;
   RECT 52.82 66.69 203.3 68.4 ;
   RECT 52.82 68.4 203.3 70.11 ;
   RECT 52.82 70.11 203.3 71.82 ;
   RECT 52.82 71.82 203.3 73.53 ;
   RECT 52.82 73.53 203.3 75.24 ;
   RECT 52.82 75.24 203.3 76.95 ;
   RECT 52.82 76.95 203.3 78.66 ;
   RECT 52.82 78.66 203.3 80.37 ;
   RECT 52.82 80.37 203.3 82.08 ;
   RECT 52.82 82.08 203.3 83.79 ;
   RECT 52.82 83.79 203.3 85.5 ;
   RECT 52.82 85.5 203.3 87.21 ;
   RECT 52.82 87.21 203.3 88.92 ;
   RECT 52.82 88.92 203.3 90.63 ;
   RECT 52.82 90.63 203.3 92.34 ;
   RECT 52.82 92.34 203.3 94.05 ;
   RECT 52.82 94.05 203.3 95.76 ;
   RECT 52.82 95.76 203.3 97.47 ;
   RECT 52.82 97.47 203.3 99.18 ;
   RECT 52.82 99.18 203.3 100.89 ;
   RECT 52.82 100.89 203.3 102.6 ;
   RECT 52.82 102.6 203.3 104.31 ;
   RECT 52.82 104.31 203.3 106.02 ;
   RECT 52.82 106.02 203.3 107.73 ;
   RECT 52.82 107.73 203.3 109.44 ;
   RECT 52.82 109.44 203.3 111.15 ;
   RECT 52.82 111.15 203.3 112.86 ;
   RECT 52.82 112.86 203.3 114.57 ;
   RECT 52.82 114.57 203.3 116.28 ;
   RECT 52.82 116.28 203.3 117.99 ;
   RECT 52.82 117.99 203.3 119.7 ;
   RECT 52.82 119.7 203.3 121.41 ;
   RECT 52.82 121.41 203.3 123.12 ;
   RECT 52.82 123.12 203.3 124.83 ;
   RECT 52.82 124.83 203.3 126.54 ;
   RECT 52.82 126.54 203.3 128.25 ;
   RECT 52.82 128.25 203.3 129.96 ;
   RECT 52.82 129.96 203.3 131.67 ;
   RECT 52.82 131.67 203.3 133.38 ;
   RECT 52.82 133.38 203.3 135.09 ;
   RECT 52.82 135.09 203.3 136.8 ;
   RECT 52.82 136.8 203.3 138.51 ;
   RECT 52.82 138.51 203.3 140.22 ;
   RECT 52.82 140.22 203.3 141.93 ;
   RECT 52.82 141.93 203.3 143.64 ;
  LAYER metal2 ;
   RECT 0.0 0.0 203.3 1.71 ;
   RECT 0.0 1.71 203.3 3.42 ;
   RECT 0.0 3.42 203.3 5.13 ;
   RECT 0.0 5.13 203.3 6.84 ;
   RECT 0.0 6.84 203.3 8.55 ;
   RECT 0.0 8.55 203.3 10.26 ;
   RECT 0.0 10.26 203.3 11.97 ;
   RECT 0.0 11.97 203.3 13.68 ;
   RECT 0.0 13.68 203.3 15.39 ;
   RECT 0.0 15.39 203.3 17.1 ;
   RECT 0.0 17.1 203.3 18.81 ;
   RECT 0.0 18.81 203.3 20.52 ;
   RECT 0.0 20.52 203.3 22.23 ;
   RECT 0.0 22.23 203.3 23.94 ;
   RECT 0.0 23.94 203.3 25.65 ;
   RECT 0.0 25.65 203.3 27.36 ;
   RECT 0.0 27.36 203.3 29.07 ;
   RECT 0.0 29.07 203.3 30.78 ;
   RECT 0.0 30.78 203.3 32.49 ;
   RECT 0.0 32.49 203.3 34.2 ;
   RECT 52.82 34.2 203.3 35.91 ;
   RECT 52.82 35.91 203.3 37.62 ;
   RECT 52.82 37.62 203.3 39.33 ;
   RECT 52.82 39.33 203.3 41.04 ;
   RECT 52.82 41.04 203.3 42.75 ;
   RECT 52.82 42.75 203.3 44.46 ;
   RECT 52.82 44.46 203.3 46.17 ;
   RECT 52.82 46.17 203.3 47.88 ;
   RECT 52.82 47.88 203.3 49.59 ;
   RECT 52.82 49.59 203.3 51.3 ;
   RECT 52.82 51.3 203.3 53.01 ;
   RECT 52.82 53.01 203.3 54.72 ;
   RECT 52.82 54.72 203.3 56.43 ;
   RECT 52.82 56.43 203.3 58.14 ;
   RECT 52.82 58.14 203.3 59.85 ;
   RECT 52.82 59.85 203.3 61.56 ;
   RECT 52.82 61.56 203.3 63.27 ;
   RECT 52.82 63.27 203.3 64.98 ;
   RECT 52.82 64.98 203.3 66.69 ;
   RECT 52.82 66.69 203.3 68.4 ;
   RECT 52.82 68.4 203.3 70.11 ;
   RECT 52.82 70.11 203.3 71.82 ;
   RECT 52.82 71.82 203.3 73.53 ;
   RECT 52.82 73.53 203.3 75.24 ;
   RECT 52.82 75.24 203.3 76.95 ;
   RECT 52.82 76.95 203.3 78.66 ;
   RECT 52.82 78.66 203.3 80.37 ;
   RECT 52.82 80.37 203.3 82.08 ;
   RECT 52.82 82.08 203.3 83.79 ;
   RECT 52.82 83.79 203.3 85.5 ;
   RECT 52.82 85.5 203.3 87.21 ;
   RECT 52.82 87.21 203.3 88.92 ;
   RECT 52.82 88.92 203.3 90.63 ;
   RECT 52.82 90.63 203.3 92.34 ;
   RECT 52.82 92.34 203.3 94.05 ;
   RECT 52.82 94.05 203.3 95.76 ;
   RECT 52.82 95.76 203.3 97.47 ;
   RECT 52.82 97.47 203.3 99.18 ;
   RECT 52.82 99.18 203.3 100.89 ;
   RECT 52.82 100.89 203.3 102.6 ;
   RECT 52.82 102.6 203.3 104.31 ;
   RECT 52.82 104.31 203.3 106.02 ;
   RECT 52.82 106.02 203.3 107.73 ;
   RECT 52.82 107.73 203.3 109.44 ;
   RECT 52.82 109.44 203.3 111.15 ;
   RECT 52.82 111.15 203.3 112.86 ;
   RECT 52.82 112.86 203.3 114.57 ;
   RECT 52.82 114.57 203.3 116.28 ;
   RECT 52.82 116.28 203.3 117.99 ;
   RECT 52.82 117.99 203.3 119.7 ;
   RECT 52.82 119.7 203.3 121.41 ;
   RECT 52.82 121.41 203.3 123.12 ;
   RECT 52.82 123.12 203.3 124.83 ;
   RECT 52.82 124.83 203.3 126.54 ;
   RECT 52.82 126.54 203.3 128.25 ;
   RECT 52.82 128.25 203.3 129.96 ;
   RECT 52.82 129.96 203.3 131.67 ;
   RECT 52.82 131.67 203.3 133.38 ;
   RECT 52.82 133.38 203.3 135.09 ;
   RECT 52.82 135.09 203.3 136.8 ;
   RECT 52.82 136.8 203.3 138.51 ;
   RECT 52.82 138.51 203.3 140.22 ;
   RECT 52.82 140.22 203.3 141.93 ;
   RECT 52.82 141.93 203.3 143.64 ;
  LAYER via2 ;
   RECT 0.0 0.0 203.3 1.71 ;
   RECT 0.0 1.71 203.3 3.42 ;
   RECT 0.0 3.42 203.3 5.13 ;
   RECT 0.0 5.13 203.3 6.84 ;
   RECT 0.0 6.84 203.3 8.55 ;
   RECT 0.0 8.55 203.3 10.26 ;
   RECT 0.0 10.26 203.3 11.97 ;
   RECT 0.0 11.97 203.3 13.68 ;
   RECT 0.0 13.68 203.3 15.39 ;
   RECT 0.0 15.39 203.3 17.1 ;
   RECT 0.0 17.1 203.3 18.81 ;
   RECT 0.0 18.81 203.3 20.52 ;
   RECT 0.0 20.52 203.3 22.23 ;
   RECT 0.0 22.23 203.3 23.94 ;
   RECT 0.0 23.94 203.3 25.65 ;
   RECT 0.0 25.65 203.3 27.36 ;
   RECT 0.0 27.36 203.3 29.07 ;
   RECT 0.0 29.07 203.3 30.78 ;
   RECT 0.0 30.78 203.3 32.49 ;
   RECT 0.0 32.49 203.3 34.2 ;
   RECT 52.82 34.2 203.3 35.91 ;
   RECT 52.82 35.91 203.3 37.62 ;
   RECT 52.82 37.62 203.3 39.33 ;
   RECT 52.82 39.33 203.3 41.04 ;
   RECT 52.82 41.04 203.3 42.75 ;
   RECT 52.82 42.75 203.3 44.46 ;
   RECT 52.82 44.46 203.3 46.17 ;
   RECT 52.82 46.17 203.3 47.88 ;
   RECT 52.82 47.88 203.3 49.59 ;
   RECT 52.82 49.59 203.3 51.3 ;
   RECT 52.82 51.3 203.3 53.01 ;
   RECT 52.82 53.01 203.3 54.72 ;
   RECT 52.82 54.72 203.3 56.43 ;
   RECT 52.82 56.43 203.3 58.14 ;
   RECT 52.82 58.14 203.3 59.85 ;
   RECT 52.82 59.85 203.3 61.56 ;
   RECT 52.82 61.56 203.3 63.27 ;
   RECT 52.82 63.27 203.3 64.98 ;
   RECT 52.82 64.98 203.3 66.69 ;
   RECT 52.82 66.69 203.3 68.4 ;
   RECT 52.82 68.4 203.3 70.11 ;
   RECT 52.82 70.11 203.3 71.82 ;
   RECT 52.82 71.82 203.3 73.53 ;
   RECT 52.82 73.53 203.3 75.24 ;
   RECT 52.82 75.24 203.3 76.95 ;
   RECT 52.82 76.95 203.3 78.66 ;
   RECT 52.82 78.66 203.3 80.37 ;
   RECT 52.82 80.37 203.3 82.08 ;
   RECT 52.82 82.08 203.3 83.79 ;
   RECT 52.82 83.79 203.3 85.5 ;
   RECT 52.82 85.5 203.3 87.21 ;
   RECT 52.82 87.21 203.3 88.92 ;
   RECT 52.82 88.92 203.3 90.63 ;
   RECT 52.82 90.63 203.3 92.34 ;
   RECT 52.82 92.34 203.3 94.05 ;
   RECT 52.82 94.05 203.3 95.76 ;
   RECT 52.82 95.76 203.3 97.47 ;
   RECT 52.82 97.47 203.3 99.18 ;
   RECT 52.82 99.18 203.3 100.89 ;
   RECT 52.82 100.89 203.3 102.6 ;
   RECT 52.82 102.6 203.3 104.31 ;
   RECT 52.82 104.31 203.3 106.02 ;
   RECT 52.82 106.02 203.3 107.73 ;
   RECT 52.82 107.73 203.3 109.44 ;
   RECT 52.82 109.44 203.3 111.15 ;
   RECT 52.82 111.15 203.3 112.86 ;
   RECT 52.82 112.86 203.3 114.57 ;
   RECT 52.82 114.57 203.3 116.28 ;
   RECT 52.82 116.28 203.3 117.99 ;
   RECT 52.82 117.99 203.3 119.7 ;
   RECT 52.82 119.7 203.3 121.41 ;
   RECT 52.82 121.41 203.3 123.12 ;
   RECT 52.82 123.12 203.3 124.83 ;
   RECT 52.82 124.83 203.3 126.54 ;
   RECT 52.82 126.54 203.3 128.25 ;
   RECT 52.82 128.25 203.3 129.96 ;
   RECT 52.82 129.96 203.3 131.67 ;
   RECT 52.82 131.67 203.3 133.38 ;
   RECT 52.82 133.38 203.3 135.09 ;
   RECT 52.82 135.09 203.3 136.8 ;
   RECT 52.82 136.8 203.3 138.51 ;
   RECT 52.82 138.51 203.3 140.22 ;
   RECT 52.82 140.22 203.3 141.93 ;
   RECT 52.82 141.93 203.3 143.64 ;
  LAYER metal3 ;
   RECT 0.0 0.0 203.3 1.71 ;
   RECT 0.0 1.71 203.3 3.42 ;
   RECT 0.0 3.42 203.3 5.13 ;
   RECT 0.0 5.13 203.3 6.84 ;
   RECT 0.0 6.84 203.3 8.55 ;
   RECT 0.0 8.55 203.3 10.26 ;
   RECT 0.0 10.26 203.3 11.97 ;
   RECT 0.0 11.97 203.3 13.68 ;
   RECT 0.0 13.68 203.3 15.39 ;
   RECT 0.0 15.39 203.3 17.1 ;
   RECT 0.0 17.1 203.3 18.81 ;
   RECT 0.0 18.81 203.3 20.52 ;
   RECT 0.0 20.52 203.3 22.23 ;
   RECT 0.0 22.23 203.3 23.94 ;
   RECT 0.0 23.94 203.3 25.65 ;
   RECT 0.0 25.65 203.3 27.36 ;
   RECT 0.0 27.36 203.3 29.07 ;
   RECT 0.0 29.07 203.3 30.78 ;
   RECT 0.0 30.78 203.3 32.49 ;
   RECT 0.0 32.49 203.3 34.2 ;
   RECT 52.82 34.2 203.3 35.91 ;
   RECT 52.82 35.91 203.3 37.62 ;
   RECT 52.82 37.62 203.3 39.33 ;
   RECT 52.82 39.33 203.3 41.04 ;
   RECT 52.82 41.04 203.3 42.75 ;
   RECT 52.82 42.75 203.3 44.46 ;
   RECT 52.82 44.46 203.3 46.17 ;
   RECT 52.82 46.17 203.3 47.88 ;
   RECT 52.82 47.88 203.3 49.59 ;
   RECT 52.82 49.59 203.3 51.3 ;
   RECT 52.82 51.3 203.3 53.01 ;
   RECT 52.82 53.01 203.3 54.72 ;
   RECT 52.82 54.72 203.3 56.43 ;
   RECT 52.82 56.43 203.3 58.14 ;
   RECT 52.82 58.14 203.3 59.85 ;
   RECT 52.82 59.85 203.3 61.56 ;
   RECT 52.82 61.56 203.3 63.27 ;
   RECT 52.82 63.27 203.3 64.98 ;
   RECT 52.82 64.98 203.3 66.69 ;
   RECT 52.82 66.69 203.3 68.4 ;
   RECT 52.82 68.4 203.3 70.11 ;
   RECT 52.82 70.11 203.3 71.82 ;
   RECT 52.82 71.82 203.3 73.53 ;
   RECT 52.82 73.53 203.3 75.24 ;
   RECT 52.82 75.24 203.3 76.95 ;
   RECT 52.82 76.95 203.3 78.66 ;
   RECT 52.82 78.66 203.3 80.37 ;
   RECT 52.82 80.37 203.3 82.08 ;
   RECT 52.82 82.08 203.3 83.79 ;
   RECT 52.82 83.79 203.3 85.5 ;
   RECT 52.82 85.5 203.3 87.21 ;
   RECT 52.82 87.21 203.3 88.92 ;
   RECT 52.82 88.92 203.3 90.63 ;
   RECT 52.82 90.63 203.3 92.34 ;
   RECT 52.82 92.34 203.3 94.05 ;
   RECT 52.82 94.05 203.3 95.76 ;
   RECT 52.82 95.76 203.3 97.47 ;
   RECT 52.82 97.47 203.3 99.18 ;
   RECT 52.82 99.18 203.3 100.89 ;
   RECT 52.82 100.89 203.3 102.6 ;
   RECT 52.82 102.6 203.3 104.31 ;
   RECT 52.82 104.31 203.3 106.02 ;
   RECT 52.82 106.02 203.3 107.73 ;
   RECT 52.82 107.73 203.3 109.44 ;
   RECT 52.82 109.44 203.3 111.15 ;
   RECT 52.82 111.15 203.3 112.86 ;
   RECT 52.82 112.86 203.3 114.57 ;
   RECT 52.82 114.57 203.3 116.28 ;
   RECT 52.82 116.28 203.3 117.99 ;
   RECT 52.82 117.99 203.3 119.7 ;
   RECT 52.82 119.7 203.3 121.41 ;
   RECT 52.82 121.41 203.3 123.12 ;
   RECT 52.82 123.12 203.3 124.83 ;
   RECT 52.82 124.83 203.3 126.54 ;
   RECT 52.82 126.54 203.3 128.25 ;
   RECT 52.82 128.25 203.3 129.96 ;
   RECT 52.82 129.96 203.3 131.67 ;
   RECT 52.82 131.67 203.3 133.38 ;
   RECT 52.82 133.38 203.3 135.09 ;
   RECT 52.82 135.09 203.3 136.8 ;
   RECT 52.82 136.8 203.3 138.51 ;
   RECT 52.82 138.51 203.3 140.22 ;
   RECT 52.82 140.22 203.3 141.93 ;
   RECT 52.82 141.93 203.3 143.64 ;
  LAYER via3 ;
   RECT 0.0 0.0 203.3 1.71 ;
   RECT 0.0 1.71 203.3 3.42 ;
   RECT 0.0 3.42 203.3 5.13 ;
   RECT 0.0 5.13 203.3 6.84 ;
   RECT 0.0 6.84 203.3 8.55 ;
   RECT 0.0 8.55 203.3 10.26 ;
   RECT 0.0 10.26 203.3 11.97 ;
   RECT 0.0 11.97 203.3 13.68 ;
   RECT 0.0 13.68 203.3 15.39 ;
   RECT 0.0 15.39 203.3 17.1 ;
   RECT 0.0 17.1 203.3 18.81 ;
   RECT 0.0 18.81 203.3 20.52 ;
   RECT 0.0 20.52 203.3 22.23 ;
   RECT 0.0 22.23 203.3 23.94 ;
   RECT 0.0 23.94 203.3 25.65 ;
   RECT 0.0 25.65 203.3 27.36 ;
   RECT 0.0 27.36 203.3 29.07 ;
   RECT 0.0 29.07 203.3 30.78 ;
   RECT 0.0 30.78 203.3 32.49 ;
   RECT 0.0 32.49 203.3 34.2 ;
   RECT 52.82 34.2 203.3 35.91 ;
   RECT 52.82 35.91 203.3 37.62 ;
   RECT 52.82 37.62 203.3 39.33 ;
   RECT 52.82 39.33 203.3 41.04 ;
   RECT 52.82 41.04 203.3 42.75 ;
   RECT 52.82 42.75 203.3 44.46 ;
   RECT 52.82 44.46 203.3 46.17 ;
   RECT 52.82 46.17 203.3 47.88 ;
   RECT 52.82 47.88 203.3 49.59 ;
   RECT 52.82 49.59 203.3 51.3 ;
   RECT 52.82 51.3 203.3 53.01 ;
   RECT 52.82 53.01 203.3 54.72 ;
   RECT 52.82 54.72 203.3 56.43 ;
   RECT 52.82 56.43 203.3 58.14 ;
   RECT 52.82 58.14 203.3 59.85 ;
   RECT 52.82 59.85 203.3 61.56 ;
   RECT 52.82 61.56 203.3 63.27 ;
   RECT 52.82 63.27 203.3 64.98 ;
   RECT 52.82 64.98 203.3 66.69 ;
   RECT 52.82 66.69 203.3 68.4 ;
   RECT 52.82 68.4 203.3 70.11 ;
   RECT 52.82 70.11 203.3 71.82 ;
   RECT 52.82 71.82 203.3 73.53 ;
   RECT 52.82 73.53 203.3 75.24 ;
   RECT 52.82 75.24 203.3 76.95 ;
   RECT 52.82 76.95 203.3 78.66 ;
   RECT 52.82 78.66 203.3 80.37 ;
   RECT 52.82 80.37 203.3 82.08 ;
   RECT 52.82 82.08 203.3 83.79 ;
   RECT 52.82 83.79 203.3 85.5 ;
   RECT 52.82 85.5 203.3 87.21 ;
   RECT 52.82 87.21 203.3 88.92 ;
   RECT 52.82 88.92 203.3 90.63 ;
   RECT 52.82 90.63 203.3 92.34 ;
   RECT 52.82 92.34 203.3 94.05 ;
   RECT 52.82 94.05 203.3 95.76 ;
   RECT 52.82 95.76 203.3 97.47 ;
   RECT 52.82 97.47 203.3 99.18 ;
   RECT 52.82 99.18 203.3 100.89 ;
   RECT 52.82 100.89 203.3 102.6 ;
   RECT 52.82 102.6 203.3 104.31 ;
   RECT 52.82 104.31 203.3 106.02 ;
   RECT 52.82 106.02 203.3 107.73 ;
   RECT 52.82 107.73 203.3 109.44 ;
   RECT 52.82 109.44 203.3 111.15 ;
   RECT 52.82 111.15 203.3 112.86 ;
   RECT 52.82 112.86 203.3 114.57 ;
   RECT 52.82 114.57 203.3 116.28 ;
   RECT 52.82 116.28 203.3 117.99 ;
   RECT 52.82 117.99 203.3 119.7 ;
   RECT 52.82 119.7 203.3 121.41 ;
   RECT 52.82 121.41 203.3 123.12 ;
   RECT 52.82 123.12 203.3 124.83 ;
   RECT 52.82 124.83 203.3 126.54 ;
   RECT 52.82 126.54 203.3 128.25 ;
   RECT 52.82 128.25 203.3 129.96 ;
   RECT 52.82 129.96 203.3 131.67 ;
   RECT 52.82 131.67 203.3 133.38 ;
   RECT 52.82 133.38 203.3 135.09 ;
   RECT 52.82 135.09 203.3 136.8 ;
   RECT 52.82 136.8 203.3 138.51 ;
   RECT 52.82 138.51 203.3 140.22 ;
   RECT 52.82 140.22 203.3 141.93 ;
   RECT 52.82 141.93 203.3 143.64 ;
  LAYER metal4 ;
   RECT 0.0 0.0 203.3 1.71 ;
   RECT 0.0 1.71 203.3 3.42 ;
   RECT 0.0 3.42 203.3 5.13 ;
   RECT 0.0 5.13 203.3 6.84 ;
   RECT 0.0 6.84 203.3 8.55 ;
   RECT 0.0 8.55 203.3 10.26 ;
   RECT 0.0 10.26 203.3 11.97 ;
   RECT 0.0 11.97 203.3 13.68 ;
   RECT 0.0 13.68 203.3 15.39 ;
   RECT 0.0 15.39 203.3 17.1 ;
   RECT 0.0 17.1 203.3 18.81 ;
   RECT 0.0 18.81 203.3 20.52 ;
   RECT 0.0 20.52 203.3 22.23 ;
   RECT 0.0 22.23 203.3 23.94 ;
   RECT 0.0 23.94 203.3 25.65 ;
   RECT 0.0 25.65 203.3 27.36 ;
   RECT 0.0 27.36 203.3 29.07 ;
   RECT 0.0 29.07 203.3 30.78 ;
   RECT 0.0 30.78 203.3 32.49 ;
   RECT 0.0 32.49 203.3 34.2 ;
   RECT 52.82 34.2 203.3 35.91 ;
   RECT 52.82 35.91 203.3 37.62 ;
   RECT 52.82 37.62 203.3 39.33 ;
   RECT 52.82 39.33 203.3 41.04 ;
   RECT 52.82 41.04 203.3 42.75 ;
   RECT 52.82 42.75 203.3 44.46 ;
   RECT 52.82 44.46 203.3 46.17 ;
   RECT 52.82 46.17 203.3 47.88 ;
   RECT 52.82 47.88 203.3 49.59 ;
   RECT 52.82 49.59 203.3 51.3 ;
   RECT 52.82 51.3 203.3 53.01 ;
   RECT 52.82 53.01 203.3 54.72 ;
   RECT 52.82 54.72 203.3 56.43 ;
   RECT 52.82 56.43 203.3 58.14 ;
   RECT 52.82 58.14 203.3 59.85 ;
   RECT 52.82 59.85 203.3 61.56 ;
   RECT 52.82 61.56 203.3 63.27 ;
   RECT 52.82 63.27 203.3 64.98 ;
   RECT 52.82 64.98 203.3 66.69 ;
   RECT 52.82 66.69 203.3 68.4 ;
   RECT 52.82 68.4 203.3 70.11 ;
   RECT 52.82 70.11 203.3 71.82 ;
   RECT 52.82 71.82 203.3 73.53 ;
   RECT 52.82 73.53 203.3 75.24 ;
   RECT 52.82 75.24 203.3 76.95 ;
   RECT 52.82 76.95 203.3 78.66 ;
   RECT 52.82 78.66 203.3 80.37 ;
   RECT 52.82 80.37 203.3 82.08 ;
   RECT 52.82 82.08 203.3 83.79 ;
   RECT 52.82 83.79 203.3 85.5 ;
   RECT 52.82 85.5 203.3 87.21 ;
   RECT 52.82 87.21 203.3 88.92 ;
   RECT 52.82 88.92 203.3 90.63 ;
   RECT 52.82 90.63 203.3 92.34 ;
   RECT 52.82 92.34 203.3 94.05 ;
   RECT 52.82 94.05 203.3 95.76 ;
   RECT 52.82 95.76 203.3 97.47 ;
   RECT 52.82 97.47 203.3 99.18 ;
   RECT 52.82 99.18 203.3 100.89 ;
   RECT 52.82 100.89 203.3 102.6 ;
   RECT 52.82 102.6 203.3 104.31 ;
   RECT 52.82 104.31 203.3 106.02 ;
   RECT 52.82 106.02 203.3 107.73 ;
   RECT 52.82 107.73 203.3 109.44 ;
   RECT 52.82 109.44 203.3 111.15 ;
   RECT 52.82 111.15 203.3 112.86 ;
   RECT 52.82 112.86 203.3 114.57 ;
   RECT 52.82 114.57 203.3 116.28 ;
   RECT 52.82 116.28 203.3 117.99 ;
   RECT 52.82 117.99 203.3 119.7 ;
   RECT 52.82 119.7 203.3 121.41 ;
   RECT 52.82 121.41 203.3 123.12 ;
   RECT 52.82 123.12 203.3 124.83 ;
   RECT 52.82 124.83 203.3 126.54 ;
   RECT 52.82 126.54 203.3 128.25 ;
   RECT 52.82 128.25 203.3 129.96 ;
   RECT 52.82 129.96 203.3 131.67 ;
   RECT 52.82 131.67 203.3 133.38 ;
   RECT 52.82 133.38 203.3 135.09 ;
   RECT 52.82 135.09 203.3 136.8 ;
   RECT 52.82 136.8 203.3 138.51 ;
   RECT 52.82 138.51 203.3 140.22 ;
   RECT 52.82 140.22 203.3 141.93 ;
   RECT 52.82 141.93 203.3 143.64 ;
 END
END block_535x756_102

MACRO block_197x180_32
 CLASS BLOCK ;
 FOREIGN block_197x180_32 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 74.86 BY 34.2 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 25.175 71.725 25.745 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 16.815 71.725 17.385 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 15.295 3.325 15.865 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 16.055 3.325 16.625 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 16.815 3.325 17.385 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 17.575 3.325 18.145 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 18.335 3.325 18.905 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 12.635 3.325 13.205 ;
  END
 END o7
 PIN o8
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 18.335 71.725 18.905 ;
  END
 END o8
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 21.375 71.725 21.945 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 70.395 21.755 70.965 22.325 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 22.135 71.725 22.705 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 70.395 22.515 70.965 23.085 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 24.415 71.725 24.985 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 70.395 24.795 70.965 25.365 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 26.695 71.725 27.265 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 27.455 71.725 28.025 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 5.035 3.325 5.605 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 16.055 71.725 16.625 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 13.775 71.725 14.345 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 12.255 71.725 12.825 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 28.975 71.725 29.545 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 25.935 71.725 26.505 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 29.735 3.325 30.305 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 17.575 71.725 18.145 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 22.895 71.725 23.465 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 4.275 71.725 4.845 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 5.035 71.725 5.605 ;
  END
 END i18
 PIN i19
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 6.935 71.725 7.505 ;
  END
 END i19
 PIN i20
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 7.695 71.725 8.265 ;
  END
 END i20
 PIN i21
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 8.835 71.725 9.405 ;
  END
 END i21
 PIN i22
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 71.155 9.595 71.725 10.165 ;
  END
 END i22
 OBS
  LAYER metal1 ;
   RECT 0 0 74.86 34.2 ;
  LAYER via1 ;
   RECT 0 0 74.86 34.2 ;
  LAYER metal2 ;
   RECT 0 0 74.86 34.2 ;
  LAYER via2 ;
   RECT 0 0 74.86 34.2 ;
  LAYER metal3 ;
   RECT 0 0 74.86 34.2 ;
  LAYER via3 ;
   RECT 0 0 74.86 34.2 ;
  LAYER metal4 ;
   RECT 0 0 74.86 34.2 ;
 END
END block_197x180_32

MACRO block_533x4428_789
 CLASS BLOCK ;
 FOREIGN block_533x4428_789 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 202.54 BY 841.32 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 834.955 26.885 835.525 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 830.775 26.885 831.345 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 794.105 26.885 794.675 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 360.715 26.885 361.285 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 356.535 26.885 357.105 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 352.545 26.885 353.115 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 348.365 26.885 348.935 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 344.375 26.885 344.945 ;
  END
 END o7
 PIN o8
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 340.195 26.885 340.765 ;
  END
 END o8
 PIN o9
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 336.205 26.885 336.775 ;
  END
 END o9
 PIN o10
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 332.025 26.885 332.595 ;
  END
 END o10
 PIN o11
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 328.035 26.885 328.605 ;
  END
 END o11
 PIN o12
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 323.855 26.885 324.425 ;
  END
 END o12
 PIN o13
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 789.925 26.885 790.495 ;
  END
 END o13
 PIN o14
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 319.865 26.885 320.435 ;
  END
 END o14
 PIN o15
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 315.685 26.885 316.255 ;
  END
 END o15
 PIN o16
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 293.455 26.885 294.025 ;
  END
 END o16
 PIN o17
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 289.275 26.885 289.845 ;
  END
 END o17
 PIN o18
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 285.285 26.885 285.855 ;
  END
 END o18
 PIN o19
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 281.105 26.885 281.675 ;
  END
 END o19
 PIN o20
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 277.115 26.885 277.685 ;
  END
 END o20
 PIN o21
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 272.935 26.885 273.505 ;
  END
 END o21
 PIN o22
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 268.945 26.885 269.515 ;
  END
 END o22
 PIN o23
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 264.765 26.885 265.335 ;
  END
 END o23
 PIN o24
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 785.935 26.885 786.505 ;
  END
 END o24
 PIN o25
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 260.775 26.885 261.345 ;
  END
 END o25
 PIN o26
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 256.595 26.885 257.165 ;
  END
 END o26
 PIN o27
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 252.605 26.885 253.175 ;
  END
 END o27
 PIN o28
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 248.425 26.885 248.995 ;
  END
 END o28
 PIN o29
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 244.435 26.885 245.005 ;
  END
 END o29
 PIN o30
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 240.255 26.885 240.825 ;
  END
 END o30
 PIN o31
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 236.265 26.885 236.835 ;
  END
 END o31
 PIN o32
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 232.085 26.885 232.655 ;
  END
 END o32
 PIN o33
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 228.095 26.885 228.665 ;
  END
 END o33
 PIN o34
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 223.915 26.885 224.485 ;
  END
 END o34
 PIN o35
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 781.755 26.885 782.325 ;
  END
 END o35
 PIN o36
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 219.925 26.885 220.495 ;
  END
 END o36
 PIN o37
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 215.745 26.885 216.315 ;
  END
 END o37
 PIN o38
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 211.755 26.885 212.325 ;
  END
 END o38
 PIN o39
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 207.575 26.885 208.145 ;
  END
 END o39
 PIN o40
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 198.455 26.885 199.025 ;
  END
 END o40
 PIN o41
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 194.275 26.885 194.845 ;
  END
 END o41
 PIN o42
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 190.285 26.885 190.855 ;
  END
 END o42
 PIN o43
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 186.105 26.885 186.675 ;
  END
 END o43
 PIN o44
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 182.115 26.885 182.685 ;
  END
 END o44
 PIN o45
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 177.935 26.885 178.505 ;
  END
 END o45
 PIN o46
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 777.765 26.885 778.335 ;
  END
 END o46
 PIN o47
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 173.945 26.885 174.515 ;
  END
 END o47
 PIN o48
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 169.765 26.885 170.335 ;
  END
 END o48
 PIN o49
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 165.775 26.885 166.345 ;
  END
 END o49
 PIN o50
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 161.595 26.885 162.165 ;
  END
 END o50
 PIN o51
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 157.605 26.885 158.175 ;
  END
 END o51
 PIN o52
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 153.425 26.885 153.995 ;
  END
 END o52
 PIN o53
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 149.435 26.885 150.005 ;
  END
 END o53
 PIN o54
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 145.255 26.885 145.825 ;
  END
 END o54
 PIN o55
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 141.265 26.885 141.835 ;
  END
 END o55
 PIN o56
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 137.085 26.885 137.655 ;
  END
 END o56
 PIN o57
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 773.585 26.885 774.155 ;
  END
 END o57
 PIN o58
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 133.095 26.885 133.665 ;
  END
 END o58
 PIN o59
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 128.915 26.885 129.485 ;
  END
 END o59
 PIN o60
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 124.925 26.885 125.495 ;
  END
 END o60
 PIN o61
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 120.745 26.885 121.315 ;
  END
 END o61
 PIN o62
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 116.755 26.885 117.325 ;
  END
 END o62
 PIN o63
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 112.575 26.885 113.145 ;
  END
 END o63
 PIN o64
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 90.345 26.885 90.915 ;
  END
 END o64
 PIN o65
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 86.165 26.885 86.735 ;
  END
 END o65
 PIN o66
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 82.175 26.885 82.745 ;
  END
 END o66
 PIN o67
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 77.995 26.885 78.565 ;
  END
 END o67
 PIN o68
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 769.595 26.885 770.165 ;
  END
 END o68
 PIN o69
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 74.005 26.885 74.575 ;
  END
 END o69
 PIN o70
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 69.825 26.885 70.395 ;
  END
 END o70
 PIN o71
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 65.835 26.885 66.405 ;
  END
 END o71
 PIN o72
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 61.655 26.885 62.225 ;
  END
 END o72
 PIN o73
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 57.665 26.885 58.235 ;
  END
 END o73
 PIN o74
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 53.485 26.885 54.055 ;
  END
 END o74
 PIN o75
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 49.495 26.885 50.065 ;
  END
 END o75
 PIN o76
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 45.315 26.885 45.885 ;
  END
 END o76
 PIN o77
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 41.325 26.885 41.895 ;
  END
 END o77
 PIN o78
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 37.145 26.885 37.715 ;
  END
 END o78
 PIN o79
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 765.415 26.885 765.985 ;
  END
 END o79
 PIN o80
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 33.155 26.885 33.725 ;
  END
 END o80
 PIN o81
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 28.975 26.885 29.545 ;
  END
 END o81
 PIN o82
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 24.985 26.885 25.555 ;
  END
 END o82
 PIN o83
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 20.805 26.885 21.375 ;
  END
 END o83
 PIN o84
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 16.815 26.885 17.385 ;
  END
 END o84
 PIN o85
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 12.635 26.885 13.205 ;
  END
 END o85
 PIN o86
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 8.645 26.885 9.215 ;
  END
 END o86
 PIN o87
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 4.465 26.885 5.035 ;
  END
 END o87
 PIN o88
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 761.425 26.885 761.995 ;
  END
 END o88
 PIN o89
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 757.245 26.885 757.815 ;
  END
 END o89
 PIN o90
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 826.785 26.885 827.355 ;
  END
 END o90
 PIN o91
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 753.255 26.885 753.825 ;
  END
 END o91
 PIN o92
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 749.075 26.885 749.645 ;
  END
 END o92
 PIN o93
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 745.085 26.885 745.655 ;
  END
 END o93
 PIN o94
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 722.665 26.885 723.235 ;
  END
 END o94
 PIN o95
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 718.675 26.885 719.245 ;
  END
 END o95
 PIN o96
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 714.495 26.885 715.065 ;
  END
 END o96
 PIN o97
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 710.505 26.885 711.075 ;
  END
 END o97
 PIN o98
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 706.325 26.885 706.895 ;
  END
 END o98
 PIN o99
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 702.335 26.885 702.905 ;
  END
 END o99
 PIN o100
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 698.155 26.885 698.725 ;
  END
 END o100
 PIN o101
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 822.605 26.885 823.175 ;
  END
 END o101
 PIN o102
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 694.165 26.885 694.735 ;
  END
 END o102
 PIN o103
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 689.985 26.885 690.555 ;
  END
 END o103
 PIN o104
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 685.995 26.885 686.565 ;
  END
 END o104
 PIN o105
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 681.815 26.885 682.385 ;
  END
 END o105
 PIN o106
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 677.825 26.885 678.395 ;
  END
 END o106
 PIN o107
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 673.645 26.885 674.215 ;
  END
 END o107
 PIN o108
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 669.655 26.885 670.225 ;
  END
 END o108
 PIN o109
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 665.475 26.885 666.045 ;
  END
 END o109
 PIN o110
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 661.485 26.885 662.055 ;
  END
 END o110
 PIN o111
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 657.305 26.885 657.875 ;
  END
 END o111
 PIN o112
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 818.615 26.885 819.185 ;
  END
 END o112
 PIN o113
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 653.315 26.885 653.885 ;
  END
 END o113
 PIN o114
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 649.135 26.885 649.705 ;
  END
 END o114
 PIN o115
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 645.145 26.885 645.715 ;
  END
 END o115
 PIN o116
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 640.965 26.885 641.535 ;
  END
 END o116
 PIN o117
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 636.975 26.885 637.545 ;
  END
 END o117
 PIN o118
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 632.795 26.885 633.365 ;
  END
 END o118
 PIN o119
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 623.675 26.885 624.245 ;
  END
 END o119
 PIN o120
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 619.495 26.885 620.065 ;
  END
 END o120
 PIN o121
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 615.505 26.885 616.075 ;
  END
 END o121
 PIN o122
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 611.325 26.885 611.895 ;
  END
 END o122
 PIN o123
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 814.435 26.885 815.005 ;
  END
 END o123
 PIN o124
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 607.335 26.885 607.905 ;
  END
 END o124
 PIN o125
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 603.155 26.885 603.725 ;
  END
 END o125
 PIN o126
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 599.165 26.885 599.735 ;
  END
 END o126
 PIN o127
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 594.985 26.885 595.555 ;
  END
 END o127
 PIN o128
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 590.995 26.885 591.565 ;
  END
 END o128
 PIN o129
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 586.815 26.885 587.385 ;
  END
 END o129
 PIN o130
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 582.825 26.885 583.395 ;
  END
 END o130
 PIN o131
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 578.645 26.885 579.215 ;
  END
 END o131
 PIN o132
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 574.655 26.885 575.225 ;
  END
 END o132
 PIN o133
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 570.475 26.885 571.045 ;
  END
 END o133
 PIN o134
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 810.445 26.885 811.015 ;
  END
 END o134
 PIN o135
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 566.485 26.885 567.055 ;
  END
 END o135
 PIN o136
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 562.305 26.885 562.875 ;
  END
 END o136
 PIN o137
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 558.315 26.885 558.885 ;
  END
 END o137
 PIN o138
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 554.135 26.885 554.705 ;
  END
 END o138
 PIN o139
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 550.145 26.885 550.715 ;
  END
 END o139
 PIN o140
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 545.965 26.885 546.535 ;
  END
 END o140
 PIN o141
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 541.975 26.885 542.545 ;
  END
 END o141
 PIN o142
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 537.795 26.885 538.365 ;
  END
 END o142
 PIN o143
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 515.565 26.885 516.135 ;
  END
 END o143
 PIN o144
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 511.385 26.885 511.955 ;
  END
 END o144
 PIN o145
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 806.265 26.885 806.835 ;
  END
 END o145
 PIN o146
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 507.395 26.885 507.965 ;
  END
 END o146
 PIN o147
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 503.215 26.885 503.785 ;
  END
 END o147
 PIN o148
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 499.225 26.885 499.795 ;
  END
 END o148
 PIN o149
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 495.045 26.885 495.615 ;
  END
 END o149
 PIN o150
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 491.055 26.885 491.625 ;
  END
 END o150
 PIN o151
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 486.875 26.885 487.445 ;
  END
 END o151
 PIN o152
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 482.885 26.885 483.455 ;
  END
 END o152
 PIN o153
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 478.705 26.885 479.275 ;
  END
 END o153
 PIN o154
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 474.715 26.885 475.285 ;
  END
 END o154
 PIN o155
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 470.535 26.885 471.105 ;
  END
 END o155
 PIN o156
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 802.275 26.885 802.845 ;
  END
 END o156
 PIN o157
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 466.545 26.885 467.115 ;
  END
 END o157
 PIN o158
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 462.365 26.885 462.935 ;
  END
 END o158
 PIN o159
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 458.375 26.885 458.945 ;
  END
 END o159
 PIN o160
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 454.195 26.885 454.765 ;
  END
 END o160
 PIN o161
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 450.205 26.885 450.775 ;
  END
 END o161
 PIN o162
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 446.025 26.885 446.595 ;
  END
 END o162
 PIN o163
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 442.035 26.885 442.605 ;
  END
 END o163
 PIN o164
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 437.855 26.885 438.425 ;
  END
 END o164
 PIN o165
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 433.865 26.885 434.435 ;
  END
 END o165
 PIN o166
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 429.685 26.885 430.255 ;
  END
 END o166
 PIN o167
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 798.095 26.885 798.665 ;
  END
 END o167
 PIN o168
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 401.565 26.885 402.135 ;
  END
 END o168
 PIN o169
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 397.385 26.885 397.955 ;
  END
 END o169
 PIN o170
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 393.395 26.885 393.965 ;
  END
 END o170
 PIN o171
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 389.215 26.885 389.785 ;
  END
 END o171
 PIN o172
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 385.225 26.885 385.795 ;
  END
 END o172
 PIN o173
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 381.045 26.885 381.615 ;
  END
 END o173
 PIN o174
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 377.055 26.885 377.625 ;
  END
 END o174
 PIN o175
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 372.875 26.885 373.445 ;
  END
 END o175
 PIN o176
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 368.885 26.885 369.455 ;
  END
 END o176
 PIN o177
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 364.705 26.885 365.275 ;
  END
 END o177
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 426.835 3.705 427.405 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 409.735 3.705 410.305 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 421.515 3.705 422.085 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 426.455 4.465 427.025 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 427.215 4.465 427.785 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 427.595 3.705 428.165 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 417.905 3.705 418.475 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 404.795 3.705 405.365 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 410.115 4.465 410.685 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 410.495 3.705 411.065 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 408.405 3.705 408.975 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 405.935 3.705 406.505 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 404.415 4.465 404.985 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 13.015 427.975 13.585 428.545 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 13.015 414.675 13.585 415.245 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 836.665 26.885 837.235 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 832.485 26.885 833.055 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 795.815 26.885 796.385 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 359.005 26.885 359.575 ;
  END
 END i18
 PIN i19
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 354.825 26.885 355.395 ;
  END
 END i19
 PIN i20
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 350.835 26.885 351.405 ;
  END
 END i20
 PIN i21
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 346.655 26.885 347.225 ;
  END
 END i21
 PIN i22
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 342.665 26.885 343.235 ;
  END
 END i22
 PIN i23
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 338.485 26.885 339.055 ;
  END
 END i23
 PIN i24
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 334.495 26.885 335.065 ;
  END
 END i24
 PIN i25
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 330.315 26.885 330.885 ;
  END
 END i25
 PIN i26
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 326.325 26.885 326.895 ;
  END
 END i26
 PIN i27
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 322.145 26.885 322.715 ;
  END
 END i27
 PIN i28
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 791.635 26.885 792.205 ;
  END
 END i28
 PIN i29
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 318.155 26.885 318.725 ;
  END
 END i29
 PIN i30
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 313.975 26.885 314.545 ;
  END
 END i30
 PIN i31
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 291.745 26.885 292.315 ;
  END
 END i31
 PIN i32
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 287.565 26.885 288.135 ;
  END
 END i32
 PIN i33
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 283.575 26.885 284.145 ;
  END
 END i33
 PIN i34
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 279.395 26.885 279.965 ;
  END
 END i34
 PIN i35
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 275.405 26.885 275.975 ;
  END
 END i35
 PIN i36
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 271.225 26.885 271.795 ;
  END
 END i36
 PIN i37
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 267.235 26.885 267.805 ;
  END
 END i37
 PIN i38
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 263.055 26.885 263.625 ;
  END
 END i38
 PIN i39
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 787.645 26.885 788.215 ;
  END
 END i39
 PIN i40
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 259.065 26.885 259.635 ;
  END
 END i40
 PIN i41
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 254.885 26.885 255.455 ;
  END
 END i41
 PIN i42
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 250.895 26.885 251.465 ;
  END
 END i42
 PIN i43
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 246.715 26.885 247.285 ;
  END
 END i43
 PIN i44
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 242.725 26.885 243.295 ;
  END
 END i44
 PIN i45
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 238.545 26.885 239.115 ;
  END
 END i45
 PIN i46
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 234.555 26.885 235.125 ;
  END
 END i46
 PIN i47
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 230.375 26.885 230.945 ;
  END
 END i47
 PIN i48
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 226.385 26.885 226.955 ;
  END
 END i48
 PIN i49
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 222.205 26.885 222.775 ;
  END
 END i49
 PIN i50
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 783.465 26.885 784.035 ;
  END
 END i50
 PIN i51
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 218.215 26.885 218.785 ;
  END
 END i51
 PIN i52
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 214.035 26.885 214.605 ;
  END
 END i52
 PIN i53
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 210.045 26.885 210.615 ;
  END
 END i53
 PIN i54
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 205.865 26.885 206.435 ;
  END
 END i54
 PIN i55
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 196.745 26.885 197.315 ;
  END
 END i55
 PIN i56
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 192.565 26.885 193.135 ;
  END
 END i56
 PIN i57
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 188.575 26.885 189.145 ;
  END
 END i57
 PIN i58
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 184.395 26.885 184.965 ;
  END
 END i58
 PIN i59
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 180.405 26.885 180.975 ;
  END
 END i59
 PIN i60
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 176.225 26.885 176.795 ;
  END
 END i60
 PIN i61
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 779.475 26.885 780.045 ;
  END
 END i61
 PIN i62
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 172.235 26.885 172.805 ;
  END
 END i62
 PIN i63
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 168.055 26.885 168.625 ;
  END
 END i63
 PIN i64
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 164.065 26.885 164.635 ;
  END
 END i64
 PIN i65
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 159.885 26.885 160.455 ;
  END
 END i65
 PIN i66
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 155.895 26.885 156.465 ;
  END
 END i66
 PIN i67
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 151.715 26.885 152.285 ;
  END
 END i67
 PIN i68
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 147.725 26.885 148.295 ;
  END
 END i68
 PIN i69
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 143.545 26.885 144.115 ;
  END
 END i69
 PIN i70
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 139.555 26.885 140.125 ;
  END
 END i70
 PIN i71
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 135.375 26.885 135.945 ;
  END
 END i71
 PIN i72
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 775.295 26.885 775.865 ;
  END
 END i72
 PIN i73
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 131.385 26.885 131.955 ;
  END
 END i73
 PIN i74
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 127.205 26.885 127.775 ;
  END
 END i74
 PIN i75
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 123.215 26.885 123.785 ;
  END
 END i75
 PIN i76
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 119.035 26.885 119.605 ;
  END
 END i76
 PIN i77
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 115.045 26.885 115.615 ;
  END
 END i77
 PIN i78
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 110.865 26.885 111.435 ;
  END
 END i78
 PIN i79
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 88.635 26.885 89.205 ;
  END
 END i79
 PIN i80
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 84.455 26.885 85.025 ;
  END
 END i80
 PIN i81
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 80.465 26.885 81.035 ;
  END
 END i81
 PIN i82
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 76.285 26.885 76.855 ;
  END
 END i82
 PIN i83
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 771.305 26.885 771.875 ;
  END
 END i83
 PIN i84
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 72.295 26.885 72.865 ;
  END
 END i84
 PIN i85
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 68.115 26.885 68.685 ;
  END
 END i85
 PIN i86
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 64.125 26.885 64.695 ;
  END
 END i86
 PIN i87
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 59.945 26.885 60.515 ;
  END
 END i87
 PIN i88
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 55.955 26.885 56.525 ;
  END
 END i88
 PIN i89
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 51.775 26.885 52.345 ;
  END
 END i89
 PIN i90
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 47.785 26.885 48.355 ;
  END
 END i90
 PIN i91
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 43.605 26.885 44.175 ;
  END
 END i91
 PIN i92
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 39.615 26.885 40.185 ;
  END
 END i92
 PIN i93
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 35.435 26.885 36.005 ;
  END
 END i93
 PIN i94
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 767.125 26.885 767.695 ;
  END
 END i94
 PIN i95
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 31.445 26.885 32.015 ;
  END
 END i95
 PIN i96
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 27.265 26.885 27.835 ;
  END
 END i96
 PIN i97
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 23.275 26.885 23.845 ;
  END
 END i97
 PIN i98
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 19.095 26.885 19.665 ;
  END
 END i98
 PIN i99
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 15.105 26.885 15.675 ;
  END
 END i99
 PIN i100
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 10.925 26.885 11.495 ;
  END
 END i100
 PIN i101
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 6.935 26.885 7.505 ;
  END
 END i101
 PIN i102
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 2.755 26.885 3.325 ;
  END
 END i102
 PIN i103
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 763.135 26.885 763.705 ;
  END
 END i103
 PIN i104
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 758.955 26.885 759.525 ;
  END
 END i104
 PIN i105
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 828.495 26.885 829.065 ;
  END
 END i105
 PIN i106
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 754.965 26.885 755.535 ;
  END
 END i106
 PIN i107
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 750.785 26.885 751.355 ;
  END
 END i107
 PIN i108
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 746.795 26.885 747.365 ;
  END
 END i108
 PIN i109
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 724.375 26.885 724.945 ;
  END
 END i109
 PIN i110
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 720.385 26.885 720.955 ;
  END
 END i110
 PIN i111
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 716.205 26.885 716.775 ;
  END
 END i111
 PIN i112
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 712.215 26.885 712.785 ;
  END
 END i112
 PIN i113
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 708.035 26.885 708.605 ;
  END
 END i113
 PIN i114
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 704.045 26.885 704.615 ;
  END
 END i114
 PIN i115
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 699.865 26.885 700.435 ;
  END
 END i115
 PIN i116
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 824.315 26.885 824.885 ;
  END
 END i116
 PIN i117
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 695.875 26.885 696.445 ;
  END
 END i117
 PIN i118
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 691.695 26.885 692.265 ;
  END
 END i118
 PIN i119
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 687.705 26.885 688.275 ;
  END
 END i119
 PIN i120
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 683.525 26.885 684.095 ;
  END
 END i120
 PIN i121
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 679.535 26.885 680.105 ;
  END
 END i121
 PIN i122
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 675.355 26.885 675.925 ;
  END
 END i122
 PIN i123
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 671.365 26.885 671.935 ;
  END
 END i123
 PIN i124
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 667.185 26.885 667.755 ;
  END
 END i124
 PIN i125
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 663.195 26.885 663.765 ;
  END
 END i125
 PIN i126
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 659.015 26.885 659.585 ;
  END
 END i126
 PIN i127
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 820.325 26.885 820.895 ;
  END
 END i127
 PIN i128
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 655.025 26.885 655.595 ;
  END
 END i128
 PIN i129
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 650.845 26.885 651.415 ;
  END
 END i129
 PIN i130
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 646.855 26.885 647.425 ;
  END
 END i130
 PIN i131
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 642.675 26.885 643.245 ;
  END
 END i131
 PIN i132
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 638.685 26.885 639.255 ;
  END
 END i132
 PIN i133
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 634.505 26.885 635.075 ;
  END
 END i133
 PIN i134
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 625.385 26.885 625.955 ;
  END
 END i134
 PIN i135
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 621.205 26.885 621.775 ;
  END
 END i135
 PIN i136
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 617.215 26.885 617.785 ;
  END
 END i136
 PIN i137
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 613.035 26.885 613.605 ;
  END
 END i137
 PIN i138
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 816.145 26.885 816.715 ;
  END
 END i138
 PIN i139
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 609.045 26.885 609.615 ;
  END
 END i139
 PIN i140
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 604.865 26.885 605.435 ;
  END
 END i140
 PIN i141
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 600.875 26.885 601.445 ;
  END
 END i141
 PIN i142
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 596.695 26.885 597.265 ;
  END
 END i142
 PIN i143
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 592.705 26.885 593.275 ;
  END
 END i143
 PIN i144
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 588.525 26.885 589.095 ;
  END
 END i144
 PIN i145
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 584.535 26.885 585.105 ;
  END
 END i145
 PIN i146
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 580.355 26.885 580.925 ;
  END
 END i146
 PIN i147
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 576.365 26.885 576.935 ;
  END
 END i147
 PIN i148
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 572.185 26.885 572.755 ;
  END
 END i148
 PIN i149
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 812.155 26.885 812.725 ;
  END
 END i149
 PIN i150
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 568.195 26.885 568.765 ;
  END
 END i150
 PIN i151
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 564.015 26.885 564.585 ;
  END
 END i151
 PIN i152
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 560.025 26.885 560.595 ;
  END
 END i152
 PIN i153
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 555.845 26.885 556.415 ;
  END
 END i153
 PIN i154
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 551.855 26.885 552.425 ;
  END
 END i154
 PIN i155
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 547.675 26.885 548.245 ;
  END
 END i155
 PIN i156
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 543.685 26.885 544.255 ;
  END
 END i156
 PIN i157
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 539.505 26.885 540.075 ;
  END
 END i157
 PIN i158
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 517.275 26.885 517.845 ;
  END
 END i158
 PIN i159
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 513.095 26.885 513.665 ;
  END
 END i159
 PIN i160
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 807.975 26.885 808.545 ;
  END
 END i160
 PIN i161
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 509.105 26.885 509.675 ;
  END
 END i161
 PIN i162
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 504.925 26.885 505.495 ;
  END
 END i162
 PIN i163
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 500.935 26.885 501.505 ;
  END
 END i163
 PIN i164
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 496.755 26.885 497.325 ;
  END
 END i164
 PIN i165
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 492.765 26.885 493.335 ;
  END
 END i165
 PIN i166
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 488.585 26.885 489.155 ;
  END
 END i166
 PIN i167
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 484.595 26.885 485.165 ;
  END
 END i167
 PIN i168
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 480.415 26.885 480.985 ;
  END
 END i168
 PIN i169
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 476.425 26.885 476.995 ;
  END
 END i169
 PIN i170
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 472.245 26.885 472.815 ;
  END
 END i170
 PIN i171
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 803.985 26.885 804.555 ;
  END
 END i171
 PIN i172
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 468.255 26.885 468.825 ;
  END
 END i172
 PIN i173
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 464.075 26.885 464.645 ;
  END
 END i173
 PIN i174
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 460.085 26.885 460.655 ;
  END
 END i174
 PIN i175
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 455.905 26.885 456.475 ;
  END
 END i175
 PIN i176
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 451.915 26.885 452.485 ;
  END
 END i176
 PIN i177
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 447.735 26.885 448.305 ;
  END
 END i177
 PIN i178
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 443.745 26.885 444.315 ;
  END
 END i178
 PIN i179
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 439.565 26.885 440.135 ;
  END
 END i179
 PIN i180
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 435.575 26.885 436.145 ;
  END
 END i180
 PIN i181
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 431.395 26.885 431.965 ;
  END
 END i181
 PIN i182
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 799.805 26.885 800.375 ;
  END
 END i182
 PIN i183
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 399.855 26.885 400.425 ;
  END
 END i183
 PIN i184
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 395.675 26.885 396.245 ;
  END
 END i184
 PIN i185
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 391.685 26.885 392.255 ;
  END
 END i185
 PIN i186
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 387.505 26.885 388.075 ;
  END
 END i186
 PIN i187
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 383.515 26.885 384.085 ;
  END
 END i187
 PIN i188
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 379.335 26.885 379.905 ;
  END
 END i188
 PIN i189
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 375.345 26.885 375.915 ;
  END
 END i189
 PIN i190
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 371.165 26.885 371.735 ;
  END
 END i190
 PIN i191
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 367.175 26.885 367.745 ;
  END
 END i191
 PIN i192
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 26.315 362.995 26.885 363.565 ;
  END
 END i192
 PIN i193
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 769.025 27.645 769.595 ;
  END
 END i193
 PIN i194
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 764.845 27.645 765.415 ;
  END
 END i194
 PIN i195
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 760.855 27.645 761.425 ;
  END
 END i195
 PIN i196
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 781.185 27.645 781.755 ;
  END
 END i196
 PIN i197
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 777.195 27.645 777.765 ;
  END
 END i197
 PIN i198
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 701.765 27.645 702.335 ;
  END
 END i198
 PIN i199
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 697.585 27.645 698.155 ;
  END
 END i199
 PIN i200
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 693.595 27.645 694.165 ;
  END
 END i200
 PIN i201
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 689.415 27.645 689.985 ;
  END
 END i201
 PIN i202
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 685.425 27.645 685.995 ;
  END
 END i202
 PIN i203
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 561.735 27.645 562.305 ;
  END
 END i203
 PIN i204
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 557.745 27.645 558.315 ;
  END
 END i204
 PIN i205
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 553.565 27.645 554.135 ;
  END
 END i205
 PIN i206
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 574.085 27.645 574.655 ;
  END
 END i206
 PIN i207
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 569.905 27.645 570.475 ;
  END
 END i207
 PIN i208
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 494.475 27.645 495.045 ;
  END
 END i208
 PIN i209
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 490.485 27.645 491.055 ;
  END
 END i209
 PIN i210
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 486.305 27.645 486.875 ;
  END
 END i210
 PIN i211
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 482.315 27.645 482.885 ;
  END
 END i211
 PIN i212
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 478.135 27.645 478.705 ;
  END
 END i212
 PIN i213
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 336.775 27.645 337.345 ;
  END
 END i213
 PIN i214
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 340.765 27.645 341.335 ;
  END
 END i214
 PIN i215
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 344.945 27.645 345.515 ;
  END
 END i215
 PIN i216
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 348.935 27.645 349.505 ;
  END
 END i216
 PIN i217
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 353.115 27.645 353.685 ;
  END
 END i217
 PIN i218
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 269.515 27.645 270.085 ;
  END
 END i218
 PIN i219
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 273.505 27.645 274.075 ;
  END
 END i219
 PIN i220
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 277.685 27.645 278.255 ;
  END
 END i220
 PIN i221
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 257.165 27.645 257.735 ;
  END
 END i221
 PIN i222
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 261.345 27.645 261.915 ;
  END
 END i222
 PIN i223
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 133.665 27.645 134.235 ;
  END
 END i223
 PIN i224
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 137.655 27.645 138.225 ;
  END
 END i224
 PIN i225
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 141.835 27.645 142.405 ;
  END
 END i225
 PIN i226
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 145.825 27.645 146.395 ;
  END
 END i226
 PIN i227
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 150.005 27.645 150.575 ;
  END
 END i227
 PIN i228
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 66.405 27.645 66.975 ;
  END
 END i228
 PIN i229
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 70.395 27.645 70.965 ;
  END
 END i229
 PIN i230
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 74.575 27.645 75.145 ;
  END
 END i230
 PIN i231
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 54.055 27.645 54.625 ;
  END
 END i231
 PIN i232
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 58.235 27.645 58.805 ;
  END
 END i232
 PIN i233
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 773.015 27.645 773.585 ;
  END
 END i233
 PIN i234
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 705.755 27.645 706.325 ;
  END
 END i234
 PIN i235
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 565.915 27.645 566.485 ;
  END
 END i235
 PIN i236
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 498.655 27.645 499.225 ;
  END
 END i236
 PIN i237
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 332.595 27.645 333.165 ;
  END
 END i237
 PIN i238
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 265.335 27.645 265.905 ;
  END
 END i238
 PIN i239
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 129.485 27.645 130.055 ;
  END
 END i239
 PIN i240
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 62.225 27.645 62.795 ;
  END
 END i240
 PIN i241
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 17.955 427.975 18.525 428.545 ;
  END
 END i241
 PIN i242
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 17.955 414.675 18.525 415.245 ;
  END
 END i242
 PIN i243
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 836.095 27.645 836.665 ;
  END
 END i243
 PIN i244
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 831.915 27.645 832.485 ;
  END
 END i244
 PIN i245
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 795.245 27.645 795.815 ;
  END
 END i245
 PIN i246
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 359.575 27.645 360.145 ;
  END
 END i246
 PIN i247
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 355.395 27.645 355.965 ;
  END
 END i247
 PIN i248
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 351.405 27.645 351.975 ;
  END
 END i248
 PIN i249
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 347.225 27.645 347.795 ;
  END
 END i249
 PIN i250
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 343.235 27.645 343.805 ;
  END
 END i250
 PIN i251
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 339.055 27.645 339.625 ;
  END
 END i251
 PIN i252
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 335.065 27.645 335.635 ;
  END
 END i252
 PIN i253
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 330.885 27.645 331.455 ;
  END
 END i253
 PIN i254
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 326.895 27.645 327.465 ;
  END
 END i254
 PIN i255
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 322.715 27.645 323.285 ;
  END
 END i255
 PIN i256
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 791.065 27.645 791.635 ;
  END
 END i256
 PIN i257
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 318.725 27.645 319.295 ;
  END
 END i257
 PIN i258
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 314.545 27.645 315.115 ;
  END
 END i258
 PIN i259
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 292.315 27.645 292.885 ;
  END
 END i259
 PIN i260
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 288.135 27.645 288.705 ;
  END
 END i260
 PIN i261
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 284.145 27.645 284.715 ;
  END
 END i261
 PIN i262
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 279.965 27.645 280.535 ;
  END
 END i262
 PIN i263
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 275.975 27.645 276.545 ;
  END
 END i263
 PIN i264
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 271.795 27.645 272.365 ;
  END
 END i264
 PIN i265
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 267.805 27.645 268.375 ;
  END
 END i265
 PIN i266
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 263.625 27.645 264.195 ;
  END
 END i266
 PIN i267
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 787.075 27.645 787.645 ;
  END
 END i267
 PIN i268
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 259.635 27.645 260.205 ;
  END
 END i268
 PIN i269
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 255.455 27.645 256.025 ;
  END
 END i269
 PIN i270
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 251.465 27.645 252.035 ;
  END
 END i270
 PIN i271
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 247.285 27.645 247.855 ;
  END
 END i271
 PIN i272
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 243.295 27.645 243.865 ;
  END
 END i272
 PIN i273
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 239.115 27.645 239.685 ;
  END
 END i273
 PIN i274
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 235.125 27.645 235.695 ;
  END
 END i274
 PIN i275
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 230.945 27.645 231.515 ;
  END
 END i275
 PIN i276
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 226.955 27.645 227.525 ;
  END
 END i276
 PIN i277
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 222.775 27.645 223.345 ;
  END
 END i277
 PIN i278
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 782.895 27.645 783.465 ;
  END
 END i278
 PIN i279
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 218.785 27.645 219.355 ;
  END
 END i279
 PIN i280
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 214.605 27.645 215.175 ;
  END
 END i280
 PIN i281
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 210.615 27.645 211.185 ;
  END
 END i281
 PIN i282
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 206.435 27.645 207.005 ;
  END
 END i282
 PIN i283
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 197.315 27.645 197.885 ;
  END
 END i283
 PIN i284
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 193.135 27.645 193.705 ;
  END
 END i284
 PIN i285
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 189.145 27.645 189.715 ;
  END
 END i285
 PIN i286
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 184.965 27.645 185.535 ;
  END
 END i286
 PIN i287
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 180.975 27.645 181.545 ;
  END
 END i287
 PIN i288
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 176.795 27.645 177.365 ;
  END
 END i288
 PIN i289
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 778.905 27.645 779.475 ;
  END
 END i289
 PIN i290
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 172.805 27.645 173.375 ;
  END
 END i290
 PIN i291
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 168.625 27.645 169.195 ;
  END
 END i291
 PIN i292
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 164.635 27.645 165.205 ;
  END
 END i292
 PIN i293
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 160.455 27.645 161.025 ;
  END
 END i293
 PIN i294
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 156.465 27.645 157.035 ;
  END
 END i294
 PIN i295
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 152.285 27.645 152.855 ;
  END
 END i295
 PIN i296
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 148.295 27.645 148.865 ;
  END
 END i296
 PIN i297
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 144.115 27.645 144.685 ;
  END
 END i297
 PIN i298
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 140.125 27.645 140.695 ;
  END
 END i298
 PIN i299
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 135.945 27.645 136.515 ;
  END
 END i299
 PIN i300
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 774.725 27.645 775.295 ;
  END
 END i300
 PIN i301
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 131.955 27.645 132.525 ;
  END
 END i301
 PIN i302
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 127.775 27.645 128.345 ;
  END
 END i302
 PIN i303
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 123.785 27.645 124.355 ;
  END
 END i303
 PIN i304
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 119.605 27.645 120.175 ;
  END
 END i304
 PIN i305
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 115.615 27.645 116.185 ;
  END
 END i305
 PIN i306
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 111.435 27.645 112.005 ;
  END
 END i306
 PIN i307
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 89.205 27.645 89.775 ;
  END
 END i307
 PIN i308
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 85.025 27.645 85.595 ;
  END
 END i308
 PIN i309
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 81.035 27.645 81.605 ;
  END
 END i309
 PIN i310
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 76.855 27.645 77.425 ;
  END
 END i310
 PIN i311
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 770.735 27.645 771.305 ;
  END
 END i311
 PIN i312
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 72.865 27.645 73.435 ;
  END
 END i312
 PIN i313
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 68.685 27.645 69.255 ;
  END
 END i313
 PIN i314
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 64.695 27.645 65.265 ;
  END
 END i314
 PIN i315
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 60.515 27.645 61.085 ;
  END
 END i315
 PIN i316
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 56.525 27.645 57.095 ;
  END
 END i316
 PIN i317
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 52.345 27.645 52.915 ;
  END
 END i317
 PIN i318
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 48.355 27.645 48.925 ;
  END
 END i318
 PIN i319
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 44.175 27.645 44.745 ;
  END
 END i319
 PIN i320
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 40.185 27.645 40.755 ;
  END
 END i320
 PIN i321
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 36.005 27.645 36.575 ;
  END
 END i321
 PIN i322
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 766.555 27.645 767.125 ;
  END
 END i322
 PIN i323
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 32.015 27.645 32.585 ;
  END
 END i323
 PIN i324
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 27.835 27.645 28.405 ;
  END
 END i324
 PIN i325
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 23.845 27.645 24.415 ;
  END
 END i325
 PIN i326
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 19.665 27.645 20.235 ;
  END
 END i326
 PIN i327
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 15.675 27.645 16.245 ;
  END
 END i327
 PIN i328
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 11.495 27.645 12.065 ;
  END
 END i328
 PIN i329
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 7.505 27.645 8.075 ;
  END
 END i329
 PIN i330
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 3.325 27.645 3.895 ;
  END
 END i330
 PIN i331
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 762.565 27.645 763.135 ;
  END
 END i331
 PIN i332
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 758.385 27.645 758.955 ;
  END
 END i332
 PIN i333
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 827.925 27.645 828.495 ;
  END
 END i333
 PIN i334
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 754.395 27.645 754.965 ;
  END
 END i334
 PIN i335
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 750.215 27.645 750.785 ;
  END
 END i335
 PIN i336
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 746.225 27.645 746.795 ;
  END
 END i336
 PIN i337
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 723.805 27.645 724.375 ;
  END
 END i337
 PIN i338
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 719.815 27.645 720.385 ;
  END
 END i338
 PIN i339
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 715.635 27.645 716.205 ;
  END
 END i339
 PIN i340
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 711.645 27.645 712.215 ;
  END
 END i340
 PIN i341
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 707.465 27.645 708.035 ;
  END
 END i341
 PIN i342
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 703.475 27.645 704.045 ;
  END
 END i342
 PIN i343
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 699.295 27.645 699.865 ;
  END
 END i343
 PIN i344
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 823.745 27.645 824.315 ;
  END
 END i344
 PIN i345
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 695.305 27.645 695.875 ;
  END
 END i345
 PIN i346
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 691.125 27.645 691.695 ;
  END
 END i346
 PIN i347
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 687.135 27.645 687.705 ;
  END
 END i347
 PIN i348
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 682.955 27.645 683.525 ;
  END
 END i348
 PIN i349
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 678.965 27.645 679.535 ;
  END
 END i349
 PIN i350
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 674.785 27.645 675.355 ;
  END
 END i350
 PIN i351
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 670.795 27.645 671.365 ;
  END
 END i351
 PIN i352
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 666.615 27.645 667.185 ;
  END
 END i352
 PIN i353
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 662.625 27.645 663.195 ;
  END
 END i353
 PIN i354
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 658.445 27.645 659.015 ;
  END
 END i354
 PIN i355
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 819.755 27.645 820.325 ;
  END
 END i355
 PIN i356
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 654.455 27.645 655.025 ;
  END
 END i356
 PIN i357
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 650.275 27.645 650.845 ;
  END
 END i357
 PIN i358
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 646.285 27.645 646.855 ;
  END
 END i358
 PIN i359
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 642.105 27.645 642.675 ;
  END
 END i359
 PIN i360
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 638.115 27.645 638.685 ;
  END
 END i360
 PIN i361
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 633.935 27.645 634.505 ;
  END
 END i361
 PIN i362
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 624.815 27.645 625.385 ;
  END
 END i362
 PIN i363
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 620.635 27.645 621.205 ;
  END
 END i363
 PIN i364
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 616.645 27.645 617.215 ;
  END
 END i364
 PIN i365
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 612.465 27.645 613.035 ;
  END
 END i365
 PIN i366
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 815.575 27.645 816.145 ;
  END
 END i366
 PIN i367
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 608.475 27.645 609.045 ;
  END
 END i367
 PIN i368
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 604.295 27.645 604.865 ;
  END
 END i368
 PIN i369
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 600.305 27.645 600.875 ;
  END
 END i369
 PIN i370
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 596.125 27.645 596.695 ;
  END
 END i370
 PIN i371
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 592.135 27.645 592.705 ;
  END
 END i371
 PIN i372
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 587.955 27.645 588.525 ;
  END
 END i372
 PIN i373
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 583.965 27.645 584.535 ;
  END
 END i373
 PIN i374
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 579.785 27.645 580.355 ;
  END
 END i374
 PIN i375
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 575.795 27.645 576.365 ;
  END
 END i375
 PIN i376
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 571.615 27.645 572.185 ;
  END
 END i376
 PIN i377
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 811.585 27.645 812.155 ;
  END
 END i377
 PIN i378
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 567.625 27.645 568.195 ;
  END
 END i378
 PIN i379
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 563.445 27.645 564.015 ;
  END
 END i379
 PIN i380
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 559.455 27.645 560.025 ;
  END
 END i380
 PIN i381
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 555.275 27.645 555.845 ;
  END
 END i381
 PIN i382
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 551.285 27.645 551.855 ;
  END
 END i382
 PIN i383
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 547.105 27.645 547.675 ;
  END
 END i383
 PIN i384
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 543.115 27.645 543.685 ;
  END
 END i384
 PIN i385
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 538.935 27.645 539.505 ;
  END
 END i385
 PIN i386
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 516.705 27.645 517.275 ;
  END
 END i386
 PIN i387
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 512.525 27.645 513.095 ;
  END
 END i387
 PIN i388
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 807.405 27.645 807.975 ;
  END
 END i388
 PIN i389
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 508.535 27.645 509.105 ;
  END
 END i389
 PIN i390
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 504.355 27.645 504.925 ;
  END
 END i390
 PIN i391
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 500.365 27.645 500.935 ;
  END
 END i391
 PIN i392
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 496.185 27.645 496.755 ;
  END
 END i392
 PIN i393
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 492.195 27.645 492.765 ;
  END
 END i393
 PIN i394
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 488.015 27.645 488.585 ;
  END
 END i394
 PIN i395
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 484.025 27.645 484.595 ;
  END
 END i395
 PIN i396
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 479.845 27.645 480.415 ;
  END
 END i396
 PIN i397
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 475.855 27.645 476.425 ;
  END
 END i397
 PIN i398
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 471.675 27.645 472.245 ;
  END
 END i398
 PIN i399
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 803.415 27.645 803.985 ;
  END
 END i399
 PIN i400
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 467.685 27.645 468.255 ;
  END
 END i400
 PIN i401
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 463.505 27.645 464.075 ;
  END
 END i401
 PIN i402
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 459.515 27.645 460.085 ;
  END
 END i402
 PIN i403
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 455.335 27.645 455.905 ;
  END
 END i403
 PIN i404
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 451.345 27.645 451.915 ;
  END
 END i404
 PIN i405
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 447.165 27.645 447.735 ;
  END
 END i405
 PIN i406
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 443.175 27.645 443.745 ;
  END
 END i406
 PIN i407
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 438.995 27.645 439.565 ;
  END
 END i407
 PIN i408
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 435.005 27.645 435.575 ;
  END
 END i408
 PIN i409
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 430.825 27.645 431.395 ;
  END
 END i409
 PIN i410
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 799.235 27.645 799.805 ;
  END
 END i410
 PIN i411
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 400.425 27.645 400.995 ;
  END
 END i411
 PIN i412
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 396.245 27.645 396.815 ;
  END
 END i412
 PIN i413
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 392.255 27.645 392.825 ;
  END
 END i413
 PIN i414
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 388.075 27.645 388.645 ;
  END
 END i414
 PIN i415
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 384.085 27.645 384.655 ;
  END
 END i415
 PIN i416
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 379.905 27.645 380.475 ;
  END
 END i416
 PIN i417
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 375.915 27.645 376.485 ;
  END
 END i417
 PIN i418
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 371.735 27.645 372.305 ;
  END
 END i418
 PIN i419
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 367.745 27.645 368.315 ;
  END
 END i419
 PIN i420
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.075 363.565 27.645 364.135 ;
  END
 END i420
 PIN i421
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.135 420.375 3.705 420.945 ;
  END
 END i421
 PIN i422
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.895 419.995 4.465 420.565 ;
  END
 END i422
 PIN i423
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 835.525 28.405 836.095 ;
  END
 END i423
 PIN i424
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 831.345 28.405 831.915 ;
  END
 END i424
 PIN i425
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 794.675 28.405 795.245 ;
  END
 END i425
 PIN i426
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 360.145 28.405 360.715 ;
  END
 END i426
 PIN i427
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 355.965 28.405 356.535 ;
  END
 END i427
 PIN i428
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 351.975 28.405 352.545 ;
  END
 END i428
 PIN i429
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 347.795 28.405 348.365 ;
  END
 END i429
 PIN i430
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 343.805 28.405 344.375 ;
  END
 END i430
 PIN i431
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 339.625 28.405 340.195 ;
  END
 END i431
 PIN i432
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 335.635 28.405 336.205 ;
  END
 END i432
 PIN i433
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 331.455 28.405 332.025 ;
  END
 END i433
 PIN i434
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 327.465 28.405 328.035 ;
  END
 END i434
 PIN i435
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 323.285 28.405 323.855 ;
  END
 END i435
 PIN i436
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 790.495 28.405 791.065 ;
  END
 END i436
 PIN i437
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 319.295 28.405 319.865 ;
  END
 END i437
 PIN i438
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 315.115 28.405 315.685 ;
  END
 END i438
 PIN i439
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 292.885 28.405 293.455 ;
  END
 END i439
 PIN i440
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 288.705 28.405 289.275 ;
  END
 END i440
 PIN i441
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 284.715 28.405 285.285 ;
  END
 END i441
 PIN i442
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 280.535 28.405 281.105 ;
  END
 END i442
 PIN i443
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 276.545 28.405 277.115 ;
  END
 END i443
 PIN i444
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 272.365 28.405 272.935 ;
  END
 END i444
 PIN i445
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 268.375 28.405 268.945 ;
  END
 END i445
 PIN i446
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 264.195 28.405 264.765 ;
  END
 END i446
 PIN i447
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 786.505 28.405 787.075 ;
  END
 END i447
 PIN i448
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 260.205 28.405 260.775 ;
  END
 END i448
 PIN i449
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 256.025 28.405 256.595 ;
  END
 END i449
 PIN i450
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 252.035 28.405 252.605 ;
  END
 END i450
 PIN i451
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 247.855 28.405 248.425 ;
  END
 END i451
 PIN i452
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 243.865 28.405 244.435 ;
  END
 END i452
 PIN i453
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 239.685 28.405 240.255 ;
  END
 END i453
 PIN i454
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 235.695 28.405 236.265 ;
  END
 END i454
 PIN i455
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 231.515 28.405 232.085 ;
  END
 END i455
 PIN i456
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 227.525 28.405 228.095 ;
  END
 END i456
 PIN i457
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 223.345 28.405 223.915 ;
  END
 END i457
 PIN i458
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 782.325 28.405 782.895 ;
  END
 END i458
 PIN i459
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 219.355 28.405 219.925 ;
  END
 END i459
 PIN i460
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 215.175 28.405 215.745 ;
  END
 END i460
 PIN i461
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 211.185 28.405 211.755 ;
  END
 END i461
 PIN i462
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 207.005 28.405 207.575 ;
  END
 END i462
 PIN i463
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 197.885 28.405 198.455 ;
  END
 END i463
 PIN i464
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 193.705 28.405 194.275 ;
  END
 END i464
 PIN i465
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 189.715 28.405 190.285 ;
  END
 END i465
 PIN i466
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 185.535 28.405 186.105 ;
  END
 END i466
 PIN i467
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 181.545 28.405 182.115 ;
  END
 END i467
 PIN i468
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 177.365 28.405 177.935 ;
  END
 END i468
 PIN i469
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 778.335 28.405 778.905 ;
  END
 END i469
 PIN i470
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 173.375 28.405 173.945 ;
  END
 END i470
 PIN i471
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 169.195 28.405 169.765 ;
  END
 END i471
 PIN i472
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 165.205 28.405 165.775 ;
  END
 END i472
 PIN i473
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 161.025 28.405 161.595 ;
  END
 END i473
 PIN i474
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 157.035 28.405 157.605 ;
  END
 END i474
 PIN i475
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 152.855 28.405 153.425 ;
  END
 END i475
 PIN i476
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 148.865 28.405 149.435 ;
  END
 END i476
 PIN i477
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 144.685 28.405 145.255 ;
  END
 END i477
 PIN i478
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 140.695 28.405 141.265 ;
  END
 END i478
 PIN i479
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 136.515 28.405 137.085 ;
  END
 END i479
 PIN i480
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 774.155 28.405 774.725 ;
  END
 END i480
 PIN i481
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 132.525 28.405 133.095 ;
  END
 END i481
 PIN i482
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 128.345 28.405 128.915 ;
  END
 END i482
 PIN i483
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 124.355 28.405 124.925 ;
  END
 END i483
 PIN i484
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 120.175 28.405 120.745 ;
  END
 END i484
 PIN i485
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 116.185 28.405 116.755 ;
  END
 END i485
 PIN i486
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 112.005 28.405 112.575 ;
  END
 END i486
 PIN i487
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 89.775 28.405 90.345 ;
  END
 END i487
 PIN i488
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 85.595 28.405 86.165 ;
  END
 END i488
 PIN i489
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 81.605 28.405 82.175 ;
  END
 END i489
 PIN i490
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 77.425 28.405 77.995 ;
  END
 END i490
 PIN i491
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 770.165 28.405 770.735 ;
  END
 END i491
 PIN i492
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 73.435 28.405 74.005 ;
  END
 END i492
 PIN i493
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 69.255 28.405 69.825 ;
  END
 END i493
 PIN i494
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 65.265 28.405 65.835 ;
  END
 END i494
 PIN i495
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 61.085 28.405 61.655 ;
  END
 END i495
 PIN i496
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 57.095 28.405 57.665 ;
  END
 END i496
 PIN i497
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 52.915 28.405 53.485 ;
  END
 END i497
 PIN i498
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 48.925 28.405 49.495 ;
  END
 END i498
 PIN i499
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 44.745 28.405 45.315 ;
  END
 END i499
 PIN i500
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 40.755 28.405 41.325 ;
  END
 END i500
 PIN i501
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 36.575 28.405 37.145 ;
  END
 END i501
 PIN i502
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 765.985 28.405 766.555 ;
  END
 END i502
 PIN i503
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 32.585 28.405 33.155 ;
  END
 END i503
 PIN i504
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 28.405 28.405 28.975 ;
  END
 END i504
 PIN i505
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 24.415 28.405 24.985 ;
  END
 END i505
 PIN i506
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 20.235 28.405 20.805 ;
  END
 END i506
 PIN i507
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 16.245 28.405 16.815 ;
  END
 END i507
 PIN i508
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 12.065 28.405 12.635 ;
  END
 END i508
 PIN i509
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 8.075 28.405 8.645 ;
  END
 END i509
 PIN i510
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 3.895 28.405 4.465 ;
  END
 END i510
 PIN i511
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 761.995 28.405 762.565 ;
  END
 END i511
 PIN i512
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 757.815 28.405 758.385 ;
  END
 END i512
 PIN i513
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 827.355 28.405 827.925 ;
  END
 END i513
 PIN i514
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 753.825 28.405 754.395 ;
  END
 END i514
 PIN i515
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 749.645 28.405 750.215 ;
  END
 END i515
 PIN i516
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 745.655 28.405 746.225 ;
  END
 END i516
 PIN i517
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 723.235 28.405 723.805 ;
  END
 END i517
 PIN i518
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 719.245 28.405 719.815 ;
  END
 END i518
 PIN i519
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 715.065 28.405 715.635 ;
  END
 END i519
 PIN i520
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 711.075 28.405 711.645 ;
  END
 END i520
 PIN i521
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 706.895 28.405 707.465 ;
  END
 END i521
 PIN i522
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 702.905 28.405 703.475 ;
  END
 END i522
 PIN i523
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 698.725 28.405 699.295 ;
  END
 END i523
 PIN i524
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 823.175 28.405 823.745 ;
  END
 END i524
 PIN i525
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 694.735 28.405 695.305 ;
  END
 END i525
 PIN i526
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 690.555 28.405 691.125 ;
  END
 END i526
 PIN i527
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 686.565 28.405 687.135 ;
  END
 END i527
 PIN i528
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 682.385 28.405 682.955 ;
  END
 END i528
 PIN i529
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 678.395 28.405 678.965 ;
  END
 END i529
 PIN i530
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 674.215 28.405 674.785 ;
  END
 END i530
 PIN i531
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 670.225 28.405 670.795 ;
  END
 END i531
 PIN i532
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 666.045 28.405 666.615 ;
  END
 END i532
 PIN i533
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 662.055 28.405 662.625 ;
  END
 END i533
 PIN i534
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 657.875 28.405 658.445 ;
  END
 END i534
 PIN i535
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 819.185 28.405 819.755 ;
  END
 END i535
 PIN i536
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 653.885 28.405 654.455 ;
  END
 END i536
 PIN i537
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 649.705 28.405 650.275 ;
  END
 END i537
 PIN i538
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 645.715 28.405 646.285 ;
  END
 END i538
 PIN i539
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 641.535 28.405 642.105 ;
  END
 END i539
 PIN i540
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 637.545 28.405 638.115 ;
  END
 END i540
 PIN i541
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 633.365 28.405 633.935 ;
  END
 END i541
 PIN i542
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 624.245 28.405 624.815 ;
  END
 END i542
 PIN i543
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 620.065 28.405 620.635 ;
  END
 END i543
 PIN i544
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 616.075 28.405 616.645 ;
  END
 END i544
 PIN i545
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 611.895 28.405 612.465 ;
  END
 END i545
 PIN i546
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 815.005 28.405 815.575 ;
  END
 END i546
 PIN i547
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 607.905 28.405 608.475 ;
  END
 END i547
 PIN i548
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 603.725 28.405 604.295 ;
  END
 END i548
 PIN i549
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 599.735 28.405 600.305 ;
  END
 END i549
 PIN i550
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 595.555 28.405 596.125 ;
  END
 END i550
 PIN i551
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 591.565 28.405 592.135 ;
  END
 END i551
 PIN i552
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 587.385 28.405 587.955 ;
  END
 END i552
 PIN i553
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 583.395 28.405 583.965 ;
  END
 END i553
 PIN i554
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 579.215 28.405 579.785 ;
  END
 END i554
 PIN i555
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 575.225 28.405 575.795 ;
  END
 END i555
 PIN i556
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 571.045 28.405 571.615 ;
  END
 END i556
 PIN i557
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 811.015 28.405 811.585 ;
  END
 END i557
 PIN i558
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 567.055 28.405 567.625 ;
  END
 END i558
 PIN i559
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 562.875 28.405 563.445 ;
  END
 END i559
 PIN i560
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 558.885 28.405 559.455 ;
  END
 END i560
 PIN i561
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 554.705 28.405 555.275 ;
  END
 END i561
 PIN i562
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 550.715 28.405 551.285 ;
  END
 END i562
 PIN i563
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 546.535 28.405 547.105 ;
  END
 END i563
 PIN i564
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 542.545 28.405 543.115 ;
  END
 END i564
 PIN i565
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 538.365 28.405 538.935 ;
  END
 END i565
 PIN i566
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 516.135 28.405 516.705 ;
  END
 END i566
 PIN i567
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 511.955 28.405 512.525 ;
  END
 END i567
 PIN i568
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 806.835 28.405 807.405 ;
  END
 END i568
 PIN i569
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 507.965 28.405 508.535 ;
  END
 END i569
 PIN i570
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 503.785 28.405 504.355 ;
  END
 END i570
 PIN i571
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 499.795 28.405 500.365 ;
  END
 END i571
 PIN i572
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 495.615 28.405 496.185 ;
  END
 END i572
 PIN i573
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 491.625 28.405 492.195 ;
  END
 END i573
 PIN i574
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 487.445 28.405 488.015 ;
  END
 END i574
 PIN i575
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 483.455 28.405 484.025 ;
  END
 END i575
 PIN i576
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 479.275 28.405 479.845 ;
  END
 END i576
 PIN i577
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 475.285 28.405 475.855 ;
  END
 END i577
 PIN i578
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 471.105 28.405 471.675 ;
  END
 END i578
 PIN i579
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 802.845 28.405 803.415 ;
  END
 END i579
 PIN i580
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 467.115 28.405 467.685 ;
  END
 END i580
 PIN i581
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 462.935 28.405 463.505 ;
  END
 END i581
 PIN i582
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 458.945 28.405 459.515 ;
  END
 END i582
 PIN i583
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 454.765 28.405 455.335 ;
  END
 END i583
 PIN i584
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 450.775 28.405 451.345 ;
  END
 END i584
 PIN i585
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 446.595 28.405 447.165 ;
  END
 END i585
 PIN i586
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 442.605 28.405 443.175 ;
  END
 END i586
 PIN i587
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 438.425 28.405 438.995 ;
  END
 END i587
 PIN i588
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 434.435 28.405 435.005 ;
  END
 END i588
 PIN i589
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 430.255 28.405 430.825 ;
  END
 END i589
 PIN i590
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 798.665 28.405 799.235 ;
  END
 END i590
 PIN i591
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 400.995 28.405 401.565 ;
  END
 END i591
 PIN i592
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 396.815 28.405 397.385 ;
  END
 END i592
 PIN i593
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 392.825 28.405 393.395 ;
  END
 END i593
 PIN i594
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 388.645 28.405 389.215 ;
  END
 END i594
 PIN i595
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 384.655 28.405 385.225 ;
  END
 END i595
 PIN i596
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 380.475 28.405 381.045 ;
  END
 END i596
 PIN i597
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 376.485 28.405 377.055 ;
  END
 END i597
 PIN i598
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 372.305 28.405 372.875 ;
  END
 END i598
 PIN i599
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 368.315 28.405 368.885 ;
  END
 END i599
 PIN i600
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 27.835 364.135 28.405 364.705 ;
  END
 END i600
 PIN i601
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 4.275 427.975 4.845 428.545 ;
  END
 END i601
 PIN i602
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 5.415 427.975 5.985 428.545 ;
  END
 END i602
 PIN i603
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 6.935 427.975 7.505 428.545 ;
  END
 END i603
 PIN i604
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 8.835 427.975 9.405 428.545 ;
  END
 END i604
 PIN i605
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.975 427.975 10.545 428.545 ;
  END
 END i605
 PIN i606
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 4.275 414.675 4.845 415.245 ;
  END
 END i606
 PIN i607
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 5.415 414.675 5.985 415.245 ;
  END
 END i607
 PIN i608
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 6.935 414.675 7.505 415.245 ;
  END
 END i608
 PIN i609
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 8.835 414.675 9.405 415.245 ;
  END
 END i609
 PIN i610
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.975 414.675 10.545 415.245 ;
  END
 END i610
 OBS
  LAYER metal1 ;
   RECT 23.18 0.0 202.54 1.71 ;
   RECT 23.18 1.71 202.54 3.42 ;
   RECT 23.18 3.42 202.54 5.13 ;
   RECT 23.18 5.13 202.54 6.84 ;
   RECT 23.18 6.84 202.54 8.55 ;
   RECT 23.18 8.55 202.54 10.26 ;
   RECT 23.18 10.26 202.54 11.97 ;
   RECT 23.18 11.97 202.54 13.68 ;
   RECT 23.18 13.68 202.54 15.39 ;
   RECT 23.18 15.39 202.54 17.1 ;
   RECT 23.18 17.1 202.54 18.81 ;
   RECT 23.18 18.81 202.54 20.52 ;
   RECT 23.18 20.52 202.54 22.23 ;
   RECT 23.18 22.23 202.54 23.94 ;
   RECT 23.18 23.94 202.54 25.65 ;
   RECT 23.18 25.65 202.54 27.36 ;
   RECT 23.18 27.36 202.54 29.07 ;
   RECT 23.18 29.07 202.54 30.78 ;
   RECT 23.18 30.78 202.54 32.49 ;
   RECT 23.18 32.49 202.54 34.2 ;
   RECT 23.18 34.2 202.54 35.91 ;
   RECT 23.18 35.91 202.54 37.62 ;
   RECT 23.18 37.62 202.54 39.33 ;
   RECT 23.18 39.33 202.54 41.04 ;
   RECT 23.18 41.04 202.54 42.75 ;
   RECT 23.18 42.75 202.54 44.46 ;
   RECT 23.18 44.46 202.54 46.17 ;
   RECT 23.18 46.17 202.54 47.88 ;
   RECT 23.18 47.88 202.54 49.59 ;
   RECT 23.18 49.59 202.54 51.3 ;
   RECT 23.18 51.3 202.54 53.01 ;
   RECT 23.18 53.01 202.54 54.72 ;
   RECT 23.18 54.72 202.54 56.43 ;
   RECT 23.18 56.43 202.54 58.14 ;
   RECT 23.18 58.14 202.54 59.85 ;
   RECT 23.18 59.85 202.54 61.56 ;
   RECT 23.18 61.56 202.54 63.27 ;
   RECT 23.18 63.27 202.54 64.98 ;
   RECT 23.18 64.98 202.54 66.69 ;
   RECT 23.18 66.69 202.54 68.4 ;
   RECT 23.18 68.4 202.54 70.11 ;
   RECT 23.18 70.11 202.54 71.82 ;
   RECT 23.18 71.82 202.54 73.53 ;
   RECT 23.18 73.53 202.54 75.24 ;
   RECT 23.18 75.24 202.54 76.95 ;
   RECT 23.18 76.95 202.54 78.66 ;
   RECT 23.18 78.66 202.54 80.37 ;
   RECT 23.18 80.37 202.54 82.08 ;
   RECT 23.18 82.08 202.54 83.79 ;
   RECT 23.18 83.79 202.54 85.5 ;
   RECT 23.18 85.5 202.54 87.21 ;
   RECT 23.18 87.21 202.54 88.92 ;
   RECT 23.18 88.92 202.54 90.63 ;
   RECT 23.18 90.63 202.54 92.34 ;
   RECT 23.18 92.34 202.54 94.05 ;
   RECT 23.18 94.05 202.54 95.76 ;
   RECT 23.18 95.76 202.54 97.47 ;
   RECT 23.18 97.47 202.54 99.18 ;
   RECT 23.18 99.18 202.54 100.89 ;
   RECT 23.18 100.89 202.54 102.6 ;
   RECT 23.18 102.6 202.54 104.31 ;
   RECT 23.18 104.31 202.54 106.02 ;
   RECT 23.18 106.02 202.54 107.73 ;
   RECT 23.18 107.73 202.54 109.44 ;
   RECT 23.18 109.44 202.54 111.15 ;
   RECT 23.18 111.15 202.54 112.86 ;
   RECT 23.18 112.86 202.54 114.57 ;
   RECT 23.18 114.57 202.54 116.28 ;
   RECT 23.18 116.28 202.54 117.99 ;
   RECT 23.18 117.99 202.54 119.7 ;
   RECT 23.18 119.7 202.54 121.41 ;
   RECT 23.18 121.41 202.54 123.12 ;
   RECT 23.18 123.12 202.54 124.83 ;
   RECT 23.18 124.83 202.54 126.54 ;
   RECT 23.18 126.54 202.54 128.25 ;
   RECT 23.18 128.25 202.54 129.96 ;
   RECT 23.18 129.96 202.54 131.67 ;
   RECT 23.18 131.67 202.54 133.38 ;
   RECT 23.18 133.38 202.54 135.09 ;
   RECT 23.18 135.09 202.54 136.8 ;
   RECT 23.18 136.8 202.54 138.51 ;
   RECT 23.18 138.51 202.54 140.22 ;
   RECT 23.18 140.22 202.54 141.93 ;
   RECT 23.18 141.93 202.54 143.64 ;
   RECT 23.18 143.64 202.54 145.35 ;
   RECT 23.18 145.35 202.54 147.06 ;
   RECT 23.18 147.06 202.54 148.77 ;
   RECT 23.18 148.77 202.54 150.48 ;
   RECT 23.18 150.48 202.54 152.19 ;
   RECT 23.18 152.19 202.54 153.9 ;
   RECT 23.18 153.9 202.54 155.61 ;
   RECT 23.18 155.61 202.54 157.32 ;
   RECT 23.18 157.32 202.54 159.03 ;
   RECT 23.18 159.03 202.54 160.74 ;
   RECT 23.18 160.74 202.54 162.45 ;
   RECT 23.18 162.45 202.54 164.16 ;
   RECT 23.18 164.16 202.54 165.87 ;
   RECT 23.18 165.87 202.54 167.58 ;
   RECT 23.18 167.58 202.54 169.29 ;
   RECT 23.18 169.29 202.54 171.0 ;
   RECT 23.18 171.0 202.54 172.71 ;
   RECT 23.18 172.71 202.54 174.42 ;
   RECT 23.18 174.42 202.54 176.13 ;
   RECT 23.18 176.13 202.54 177.84 ;
   RECT 23.18 177.84 202.54 179.55 ;
   RECT 23.18 179.55 202.54 181.26 ;
   RECT 23.18 181.26 202.54 182.97 ;
   RECT 23.18 182.97 202.54 184.68 ;
   RECT 23.18 184.68 202.54 186.39 ;
   RECT 23.18 186.39 202.54 188.1 ;
   RECT 23.18 188.1 202.54 189.81 ;
   RECT 23.18 189.81 202.54 191.52 ;
   RECT 23.18 191.52 202.54 193.23 ;
   RECT 23.18 193.23 202.54 194.94 ;
   RECT 23.18 194.94 202.54 196.65 ;
   RECT 23.18 196.65 202.54 198.36 ;
   RECT 23.18 198.36 202.54 200.07 ;
   RECT 23.18 200.07 202.54 201.78 ;
   RECT 23.18 201.78 202.54 203.49 ;
   RECT 23.18 203.49 202.54 205.2 ;
   RECT 23.18 205.2 202.54 206.91 ;
   RECT 23.18 206.91 202.54 208.62 ;
   RECT 23.18 208.62 202.54 210.33 ;
   RECT 23.18 210.33 202.54 212.04 ;
   RECT 23.18 212.04 202.54 213.75 ;
   RECT 23.18 213.75 202.54 215.46 ;
   RECT 23.18 215.46 202.54 217.17 ;
   RECT 23.18 217.17 202.54 218.88 ;
   RECT 23.18 218.88 202.54 220.59 ;
   RECT 23.18 220.59 202.54 222.3 ;
   RECT 23.18 222.3 202.54 224.01 ;
   RECT 23.18 224.01 202.54 225.72 ;
   RECT 23.18 225.72 202.54 227.43 ;
   RECT 23.18 227.43 202.54 229.14 ;
   RECT 23.18 229.14 202.54 230.85 ;
   RECT 23.18 230.85 202.54 232.56 ;
   RECT 23.18 232.56 202.54 234.27 ;
   RECT 23.18 234.27 202.54 235.98 ;
   RECT 23.18 235.98 202.54 237.69 ;
   RECT 23.18 237.69 202.54 239.4 ;
   RECT 23.18 239.4 202.54 241.11 ;
   RECT 23.18 241.11 202.54 242.82 ;
   RECT 23.18 242.82 202.54 244.53 ;
   RECT 23.18 244.53 202.54 246.24 ;
   RECT 23.18 246.24 202.54 247.95 ;
   RECT 23.18 247.95 202.54 249.66 ;
   RECT 23.18 249.66 202.54 251.37 ;
   RECT 23.18 251.37 202.54 253.08 ;
   RECT 23.18 253.08 202.54 254.79 ;
   RECT 23.18 254.79 202.54 256.5 ;
   RECT 23.18 256.5 202.54 258.21 ;
   RECT 23.18 258.21 202.54 259.92 ;
   RECT 23.18 259.92 202.54 261.63 ;
   RECT 23.18 261.63 202.54 263.34 ;
   RECT 23.18 263.34 202.54 265.05 ;
   RECT 23.18 265.05 202.54 266.76 ;
   RECT 23.18 266.76 202.54 268.47 ;
   RECT 23.18 268.47 202.54 270.18 ;
   RECT 23.18 270.18 202.54 271.89 ;
   RECT 23.18 271.89 202.54 273.6 ;
   RECT 23.18 273.6 202.54 275.31 ;
   RECT 23.18 275.31 202.54 277.02 ;
   RECT 23.18 277.02 202.54 278.73 ;
   RECT 23.18 278.73 202.54 280.44 ;
   RECT 23.18 280.44 202.54 282.15 ;
   RECT 23.18 282.15 202.54 283.86 ;
   RECT 23.18 283.86 202.54 285.57 ;
   RECT 23.18 285.57 202.54 287.28 ;
   RECT 23.18 287.28 202.54 288.99 ;
   RECT 23.18 288.99 202.54 290.7 ;
   RECT 23.18 290.7 202.54 292.41 ;
   RECT 23.18 292.41 202.54 294.12 ;
   RECT 23.18 294.12 202.54 295.83 ;
   RECT 23.18 295.83 202.54 297.54 ;
   RECT 23.18 297.54 202.54 299.25 ;
   RECT 23.18 299.25 202.54 300.96 ;
   RECT 23.18 300.96 202.54 302.67 ;
   RECT 23.18 302.67 202.54 304.38 ;
   RECT 23.18 304.38 202.54 306.09 ;
   RECT 23.18 306.09 202.54 307.8 ;
   RECT 23.18 307.8 202.54 309.51 ;
   RECT 23.18 309.51 202.54 311.22 ;
   RECT 23.18 311.22 202.54 312.93 ;
   RECT 23.18 312.93 202.54 314.64 ;
   RECT 23.18 314.64 202.54 316.35 ;
   RECT 23.18 316.35 202.54 318.06 ;
   RECT 23.18 318.06 202.54 319.77 ;
   RECT 23.18 319.77 202.54 321.48 ;
   RECT 23.18 321.48 202.54 323.19 ;
   RECT 23.18 323.19 202.54 324.9 ;
   RECT 23.18 324.9 202.54 326.61 ;
   RECT 23.18 326.61 202.54 328.32 ;
   RECT 23.18 328.32 202.54 330.03 ;
   RECT 23.18 330.03 202.54 331.74 ;
   RECT 23.18 331.74 202.54 333.45 ;
   RECT 23.18 333.45 202.54 335.16 ;
   RECT 23.18 335.16 202.54 336.87 ;
   RECT 23.18 336.87 202.54 338.58 ;
   RECT 23.18 338.58 202.54 340.29 ;
   RECT 23.18 340.29 202.54 342.0 ;
   RECT 23.18 342.0 202.54 343.71 ;
   RECT 23.18 343.71 202.54 345.42 ;
   RECT 23.18 345.42 202.54 347.13 ;
   RECT 23.18 347.13 202.54 348.84 ;
   RECT 23.18 348.84 202.54 350.55 ;
   RECT 23.18 350.55 202.54 352.26 ;
   RECT 23.18 352.26 202.54 353.97 ;
   RECT 23.18 353.97 202.54 355.68 ;
   RECT 23.18 355.68 202.54 357.39 ;
   RECT 23.18 357.39 202.54 359.1 ;
   RECT 23.18 359.1 202.54 360.81 ;
   RECT 23.18 360.81 202.54 362.52 ;
   RECT 23.18 362.52 202.54 364.23 ;
   RECT 23.18 364.23 202.54 365.94 ;
   RECT 23.18 365.94 202.54 367.65 ;
   RECT 23.18 367.65 202.54 369.36 ;
   RECT 23.18 369.36 202.54 371.07 ;
   RECT 23.18 371.07 202.54 372.78 ;
   RECT 23.18 372.78 202.54 374.49 ;
   RECT 23.18 374.49 202.54 376.2 ;
   RECT 23.18 376.2 202.54 377.91 ;
   RECT 23.18 377.91 202.54 379.62 ;
   RECT 23.18 379.62 202.54 381.33 ;
   RECT 23.18 381.33 202.54 383.04 ;
   RECT 23.18 383.04 202.54 384.75 ;
   RECT 23.18 384.75 202.54 386.46 ;
   RECT 23.18 386.46 202.54 388.17 ;
   RECT 23.18 388.17 202.54 389.88 ;
   RECT 23.18 389.88 202.54 391.59 ;
   RECT 23.18 391.59 202.54 393.3 ;
   RECT 23.18 393.3 202.54 395.01 ;
   RECT 23.18 395.01 202.54 396.72 ;
   RECT 23.18 396.72 202.54 398.43 ;
   RECT 23.18 398.43 202.54 400.14 ;
   RECT 23.18 400.14 202.54 401.85 ;
   RECT 0.0 401.85 202.54 403.56 ;
   RECT 0.0 403.56 202.54 405.27 ;
   RECT 0.0 405.27 202.54 406.98 ;
   RECT 0.0 406.98 202.54 408.69 ;
   RECT 0.0 408.69 202.54 410.4 ;
   RECT 0.0 410.4 202.54 412.11 ;
   RECT 0.0 412.11 202.54 413.82 ;
   RECT 0.0 413.82 202.54 415.53 ;
   RECT 0.0 415.53 202.54 417.24 ;
   RECT 0.0 417.24 202.54 418.95 ;
   RECT 0.0 418.95 202.54 420.66 ;
   RECT 0.0 420.66 202.54 422.37 ;
   RECT 0.0 422.37 202.54 424.08 ;
   RECT 0.0 424.08 202.54 425.79 ;
   RECT 0.0 425.79 202.54 427.5 ;
   RECT 0.0 427.5 202.54 429.21 ;
   RECT 0.0 429.21 202.54 430.92 ;
   RECT 23.18 430.92 202.54 432.63 ;
   RECT 23.18 432.63 202.54 434.34 ;
   RECT 23.18 434.34 202.54 436.05 ;
   RECT 23.18 436.05 202.54 437.76 ;
   RECT 23.18 437.76 202.54 439.47 ;
   RECT 23.18 439.47 202.54 441.18 ;
   RECT 23.18 441.18 202.54 442.89 ;
   RECT 23.18 442.89 202.54 444.6 ;
   RECT 23.18 444.6 202.54 446.31 ;
   RECT 23.18 446.31 202.54 448.02 ;
   RECT 23.18 448.02 202.54 449.73 ;
   RECT 23.18 449.73 202.54 451.44 ;
   RECT 23.18 451.44 202.54 453.15 ;
   RECT 23.18 453.15 202.54 454.86 ;
   RECT 23.18 454.86 202.54 456.57 ;
   RECT 23.18 456.57 202.54 458.28 ;
   RECT 23.18 458.28 202.54 459.99 ;
   RECT 23.18 459.99 202.54 461.7 ;
   RECT 23.18 461.7 202.54 463.41 ;
   RECT 23.18 463.41 202.54 465.12 ;
   RECT 23.18 465.12 202.54 466.83 ;
   RECT 23.18 466.83 202.54 468.54 ;
   RECT 23.18 468.54 202.54 470.25 ;
   RECT 23.18 470.25 202.54 471.96 ;
   RECT 23.18 471.96 202.54 473.67 ;
   RECT 23.18 473.67 202.54 475.38 ;
   RECT 23.18 475.38 202.54 477.09 ;
   RECT 23.18 477.09 202.54 478.8 ;
   RECT 23.18 478.8 202.54 480.51 ;
   RECT 23.18 480.51 202.54 482.22 ;
   RECT 23.18 482.22 202.54 483.93 ;
   RECT 23.18 483.93 202.54 485.64 ;
   RECT 23.18 485.64 202.54 487.35 ;
   RECT 23.18 487.35 202.54 489.06 ;
   RECT 23.18 489.06 202.54 490.77 ;
   RECT 23.18 490.77 202.54 492.48 ;
   RECT 23.18 492.48 202.54 494.19 ;
   RECT 23.18 494.19 202.54 495.9 ;
   RECT 23.18 495.9 202.54 497.61 ;
   RECT 23.18 497.61 202.54 499.32 ;
   RECT 23.18 499.32 202.54 501.03 ;
   RECT 23.18 501.03 202.54 502.74 ;
   RECT 23.18 502.74 202.54 504.45 ;
   RECT 23.18 504.45 202.54 506.16 ;
   RECT 23.18 506.16 202.54 507.87 ;
   RECT 23.18 507.87 202.54 509.58 ;
   RECT 23.18 509.58 202.54 511.29 ;
   RECT 23.18 511.29 202.54 513.0 ;
   RECT 23.18 513.0 202.54 514.71 ;
   RECT 23.18 514.71 202.54 516.42 ;
   RECT 23.18 516.42 202.54 518.13 ;
   RECT 23.18 518.13 202.54 519.84 ;
   RECT 23.18 519.84 202.54 521.55 ;
   RECT 23.18 521.55 202.54 523.26 ;
   RECT 23.18 523.26 202.54 524.97 ;
   RECT 23.18 524.97 202.54 526.68 ;
   RECT 23.18 526.68 202.54 528.39 ;
   RECT 23.18 528.39 202.54 530.1 ;
   RECT 23.18 530.1 202.54 531.81 ;
   RECT 23.18 531.81 202.54 533.52 ;
   RECT 23.18 533.52 202.54 535.23 ;
   RECT 23.18 535.23 202.54 536.94 ;
   RECT 23.18 536.94 202.54 538.65 ;
   RECT 23.18 538.65 202.54 540.36 ;
   RECT 23.18 540.36 202.54 542.07 ;
   RECT 23.18 542.07 202.54 543.78 ;
   RECT 23.18 543.78 202.54 545.49 ;
   RECT 23.18 545.49 202.54 547.2 ;
   RECT 23.18 547.2 202.54 548.91 ;
   RECT 23.18 548.91 202.54 550.62 ;
   RECT 23.18 550.62 202.54 552.33 ;
   RECT 23.18 552.33 202.54 554.04 ;
   RECT 23.18 554.04 202.54 555.75 ;
   RECT 23.18 555.75 202.54 557.46 ;
   RECT 23.18 557.46 202.54 559.17 ;
   RECT 23.18 559.17 202.54 560.88 ;
   RECT 23.18 560.88 202.54 562.59 ;
   RECT 23.18 562.59 202.54 564.3 ;
   RECT 23.18 564.3 202.54 566.01 ;
   RECT 23.18 566.01 202.54 567.72 ;
   RECT 23.18 567.72 202.54 569.43 ;
   RECT 23.18 569.43 202.54 571.14 ;
   RECT 23.18 571.14 202.54 572.85 ;
   RECT 23.18 572.85 202.54 574.56 ;
   RECT 23.18 574.56 202.54 576.27 ;
   RECT 23.18 576.27 202.54 577.98 ;
   RECT 23.18 577.98 202.54 579.69 ;
   RECT 23.18 579.69 202.54 581.4 ;
   RECT 23.18 581.4 202.54 583.11 ;
   RECT 23.18 583.11 202.54 584.82 ;
   RECT 23.18 584.82 202.54 586.53 ;
   RECT 23.18 586.53 202.54 588.24 ;
   RECT 23.18 588.24 202.54 589.95 ;
   RECT 23.18 589.95 202.54 591.66 ;
   RECT 23.18 591.66 202.54 593.37 ;
   RECT 23.18 593.37 202.54 595.08 ;
   RECT 23.18 595.08 202.54 596.79 ;
   RECT 23.18 596.79 202.54 598.5 ;
   RECT 23.18 598.5 202.54 600.21 ;
   RECT 23.18 600.21 202.54 601.92 ;
   RECT 23.18 601.92 202.54 603.63 ;
   RECT 23.18 603.63 202.54 605.34 ;
   RECT 23.18 605.34 202.54 607.05 ;
   RECT 23.18 607.05 202.54 608.76 ;
   RECT 23.18 608.76 202.54 610.47 ;
   RECT 23.18 610.47 202.54 612.18 ;
   RECT 23.18 612.18 202.54 613.89 ;
   RECT 23.18 613.89 202.54 615.6 ;
   RECT 23.18 615.6 202.54 617.31 ;
   RECT 23.18 617.31 202.54 619.02 ;
   RECT 23.18 619.02 202.54 620.73 ;
   RECT 23.18 620.73 202.54 622.44 ;
   RECT 23.18 622.44 202.54 624.15 ;
   RECT 23.18 624.15 202.54 625.86 ;
   RECT 23.18 625.86 202.54 627.57 ;
   RECT 23.18 627.57 202.54 629.28 ;
   RECT 23.18 629.28 202.54 630.99 ;
   RECT 23.18 630.99 202.54 632.7 ;
   RECT 23.18 632.7 202.54 634.41 ;
   RECT 23.18 634.41 202.54 636.12 ;
   RECT 23.18 636.12 202.54 637.83 ;
   RECT 23.18 637.83 202.54 639.54 ;
   RECT 23.18 639.54 202.54 641.25 ;
   RECT 23.18 641.25 202.54 642.96 ;
   RECT 23.18 642.96 202.54 644.67 ;
   RECT 23.18 644.67 202.54 646.38 ;
   RECT 23.18 646.38 202.54 648.09 ;
   RECT 23.18 648.09 202.54 649.8 ;
   RECT 23.18 649.8 202.54 651.51 ;
   RECT 23.18 651.51 202.54 653.22 ;
   RECT 23.18 653.22 202.54 654.93 ;
   RECT 23.18 654.93 202.54 656.64 ;
   RECT 23.18 656.64 202.54 658.35 ;
   RECT 23.18 658.35 202.54 660.06 ;
   RECT 23.18 660.06 202.54 661.77 ;
   RECT 23.18 661.77 202.54 663.48 ;
   RECT 23.18 663.48 202.54 665.19 ;
   RECT 23.18 665.19 202.54 666.9 ;
   RECT 23.18 666.9 202.54 668.61 ;
   RECT 23.18 668.61 202.54 670.32 ;
   RECT 23.18 670.32 202.54 672.03 ;
   RECT 23.18 672.03 202.54 673.74 ;
   RECT 23.18 673.74 202.54 675.45 ;
   RECT 23.18 675.45 202.54 677.16 ;
   RECT 23.18 677.16 202.54 678.87 ;
   RECT 23.18 678.87 202.54 680.58 ;
   RECT 23.18 680.58 202.54 682.29 ;
   RECT 23.18 682.29 202.54 684.0 ;
   RECT 23.18 684.0 202.54 685.71 ;
   RECT 23.18 685.71 202.54 687.42 ;
   RECT 23.18 687.42 202.54 689.13 ;
   RECT 23.18 689.13 202.54 690.84 ;
   RECT 23.18 690.84 202.54 692.55 ;
   RECT 23.18 692.55 202.54 694.26 ;
   RECT 23.18 694.26 202.54 695.97 ;
   RECT 23.18 695.97 202.54 697.68 ;
   RECT 23.18 697.68 202.54 699.39 ;
   RECT 23.18 699.39 202.54 701.1 ;
   RECT 23.18 701.1 202.54 702.81 ;
   RECT 23.18 702.81 202.54 704.52 ;
   RECT 23.18 704.52 202.54 706.23 ;
   RECT 23.18 706.23 202.54 707.94 ;
   RECT 23.18 707.94 202.54 709.65 ;
   RECT 23.18 709.65 202.54 711.36 ;
   RECT 23.18 711.36 202.54 713.07 ;
   RECT 23.18 713.07 202.54 714.78 ;
   RECT 23.18 714.78 202.54 716.49 ;
   RECT 23.18 716.49 202.54 718.2 ;
   RECT 23.18 718.2 202.54 719.91 ;
   RECT 23.18 719.91 202.54 721.62 ;
   RECT 23.18 721.62 202.54 723.33 ;
   RECT 23.18 723.33 202.54 725.04 ;
   RECT 23.18 725.04 202.54 726.75 ;
   RECT 23.18 726.75 202.54 728.46 ;
   RECT 23.18 728.46 202.54 730.17 ;
   RECT 23.18 730.17 202.54 731.88 ;
   RECT 23.18 731.88 202.54 733.59 ;
   RECT 23.18 733.59 202.54 735.3 ;
   RECT 23.18 735.3 202.54 737.01 ;
   RECT 23.18 737.01 202.54 738.72 ;
   RECT 23.18 738.72 202.54 740.43 ;
   RECT 23.18 740.43 202.54 742.14 ;
   RECT 23.18 742.14 202.54 743.85 ;
   RECT 23.18 743.85 202.54 745.56 ;
   RECT 23.18 745.56 202.54 747.27 ;
   RECT 23.18 747.27 202.54 748.98 ;
   RECT 23.18 748.98 202.54 750.69 ;
   RECT 23.18 750.69 202.54 752.4 ;
   RECT 23.18 752.4 202.54 754.11 ;
   RECT 23.18 754.11 202.54 755.82 ;
   RECT 23.18 755.82 202.54 757.53 ;
   RECT 23.18 757.53 202.54 759.24 ;
   RECT 23.18 759.24 202.54 760.95 ;
   RECT 23.18 760.95 202.54 762.66 ;
   RECT 23.18 762.66 202.54 764.37 ;
   RECT 23.18 764.37 202.54 766.08 ;
   RECT 23.18 766.08 202.54 767.79 ;
   RECT 23.18 767.79 202.54 769.5 ;
   RECT 23.18 769.5 202.54 771.21 ;
   RECT 23.18 771.21 202.54 772.92 ;
   RECT 23.18 772.92 202.54 774.63 ;
   RECT 23.18 774.63 202.54 776.34 ;
   RECT 23.18 776.34 202.54 778.05 ;
   RECT 23.18 778.05 202.54 779.76 ;
   RECT 23.18 779.76 202.54 781.47 ;
   RECT 23.18 781.47 202.54 783.18 ;
   RECT 23.18 783.18 202.54 784.89 ;
   RECT 23.18 784.89 202.54 786.6 ;
   RECT 23.18 786.6 202.54 788.31 ;
   RECT 23.18 788.31 202.54 790.02 ;
   RECT 23.18 790.02 202.54 791.73 ;
   RECT 23.18 791.73 202.54 793.44 ;
   RECT 23.18 793.44 202.54 795.15 ;
   RECT 23.18 795.15 202.54 796.86 ;
   RECT 23.18 796.86 202.54 798.57 ;
   RECT 23.18 798.57 202.54 800.28 ;
   RECT 23.18 800.28 202.54 801.99 ;
   RECT 23.18 801.99 202.54 803.7 ;
   RECT 23.18 803.7 202.54 805.41 ;
   RECT 23.18 805.41 202.54 807.12 ;
   RECT 23.18 807.12 202.54 808.83 ;
   RECT 23.18 808.83 202.54 810.54 ;
   RECT 23.18 810.54 202.54 812.25 ;
   RECT 23.18 812.25 202.54 813.96 ;
   RECT 23.18 813.96 202.54 815.67 ;
   RECT 23.18 815.67 202.54 817.38 ;
   RECT 23.18 817.38 202.54 819.09 ;
   RECT 23.18 819.09 202.54 820.8 ;
   RECT 23.18 820.8 202.54 822.51 ;
   RECT 23.18 822.51 202.54 824.22 ;
   RECT 23.18 824.22 202.54 825.93 ;
   RECT 23.18 825.93 202.54 827.64 ;
   RECT 23.18 827.64 202.54 829.35 ;
   RECT 23.18 829.35 202.54 831.06 ;
   RECT 23.18 831.06 202.54 832.77 ;
   RECT 23.18 832.77 202.54 834.48 ;
   RECT 23.18 834.48 202.54 836.19 ;
   RECT 23.18 836.19 202.54 837.9 ;
   RECT 23.18 837.9 202.54 839.61 ;
   RECT 23.18 839.61 202.54 841.32 ;
  LAYER via1 ;
   RECT 23.18 0.0 202.54 1.71 ;
   RECT 23.18 1.71 202.54 3.42 ;
   RECT 23.18 3.42 202.54 5.13 ;
   RECT 23.18 5.13 202.54 6.84 ;
   RECT 23.18 6.84 202.54 8.55 ;
   RECT 23.18 8.55 202.54 10.26 ;
   RECT 23.18 10.26 202.54 11.97 ;
   RECT 23.18 11.97 202.54 13.68 ;
   RECT 23.18 13.68 202.54 15.39 ;
   RECT 23.18 15.39 202.54 17.1 ;
   RECT 23.18 17.1 202.54 18.81 ;
   RECT 23.18 18.81 202.54 20.52 ;
   RECT 23.18 20.52 202.54 22.23 ;
   RECT 23.18 22.23 202.54 23.94 ;
   RECT 23.18 23.94 202.54 25.65 ;
   RECT 23.18 25.65 202.54 27.36 ;
   RECT 23.18 27.36 202.54 29.07 ;
   RECT 23.18 29.07 202.54 30.78 ;
   RECT 23.18 30.78 202.54 32.49 ;
   RECT 23.18 32.49 202.54 34.2 ;
   RECT 23.18 34.2 202.54 35.91 ;
   RECT 23.18 35.91 202.54 37.62 ;
   RECT 23.18 37.62 202.54 39.33 ;
   RECT 23.18 39.33 202.54 41.04 ;
   RECT 23.18 41.04 202.54 42.75 ;
   RECT 23.18 42.75 202.54 44.46 ;
   RECT 23.18 44.46 202.54 46.17 ;
   RECT 23.18 46.17 202.54 47.88 ;
   RECT 23.18 47.88 202.54 49.59 ;
   RECT 23.18 49.59 202.54 51.3 ;
   RECT 23.18 51.3 202.54 53.01 ;
   RECT 23.18 53.01 202.54 54.72 ;
   RECT 23.18 54.72 202.54 56.43 ;
   RECT 23.18 56.43 202.54 58.14 ;
   RECT 23.18 58.14 202.54 59.85 ;
   RECT 23.18 59.85 202.54 61.56 ;
   RECT 23.18 61.56 202.54 63.27 ;
   RECT 23.18 63.27 202.54 64.98 ;
   RECT 23.18 64.98 202.54 66.69 ;
   RECT 23.18 66.69 202.54 68.4 ;
   RECT 23.18 68.4 202.54 70.11 ;
   RECT 23.18 70.11 202.54 71.82 ;
   RECT 23.18 71.82 202.54 73.53 ;
   RECT 23.18 73.53 202.54 75.24 ;
   RECT 23.18 75.24 202.54 76.95 ;
   RECT 23.18 76.95 202.54 78.66 ;
   RECT 23.18 78.66 202.54 80.37 ;
   RECT 23.18 80.37 202.54 82.08 ;
   RECT 23.18 82.08 202.54 83.79 ;
   RECT 23.18 83.79 202.54 85.5 ;
   RECT 23.18 85.5 202.54 87.21 ;
   RECT 23.18 87.21 202.54 88.92 ;
   RECT 23.18 88.92 202.54 90.63 ;
   RECT 23.18 90.63 202.54 92.34 ;
   RECT 23.18 92.34 202.54 94.05 ;
   RECT 23.18 94.05 202.54 95.76 ;
   RECT 23.18 95.76 202.54 97.47 ;
   RECT 23.18 97.47 202.54 99.18 ;
   RECT 23.18 99.18 202.54 100.89 ;
   RECT 23.18 100.89 202.54 102.6 ;
   RECT 23.18 102.6 202.54 104.31 ;
   RECT 23.18 104.31 202.54 106.02 ;
   RECT 23.18 106.02 202.54 107.73 ;
   RECT 23.18 107.73 202.54 109.44 ;
   RECT 23.18 109.44 202.54 111.15 ;
   RECT 23.18 111.15 202.54 112.86 ;
   RECT 23.18 112.86 202.54 114.57 ;
   RECT 23.18 114.57 202.54 116.28 ;
   RECT 23.18 116.28 202.54 117.99 ;
   RECT 23.18 117.99 202.54 119.7 ;
   RECT 23.18 119.7 202.54 121.41 ;
   RECT 23.18 121.41 202.54 123.12 ;
   RECT 23.18 123.12 202.54 124.83 ;
   RECT 23.18 124.83 202.54 126.54 ;
   RECT 23.18 126.54 202.54 128.25 ;
   RECT 23.18 128.25 202.54 129.96 ;
   RECT 23.18 129.96 202.54 131.67 ;
   RECT 23.18 131.67 202.54 133.38 ;
   RECT 23.18 133.38 202.54 135.09 ;
   RECT 23.18 135.09 202.54 136.8 ;
   RECT 23.18 136.8 202.54 138.51 ;
   RECT 23.18 138.51 202.54 140.22 ;
   RECT 23.18 140.22 202.54 141.93 ;
   RECT 23.18 141.93 202.54 143.64 ;
   RECT 23.18 143.64 202.54 145.35 ;
   RECT 23.18 145.35 202.54 147.06 ;
   RECT 23.18 147.06 202.54 148.77 ;
   RECT 23.18 148.77 202.54 150.48 ;
   RECT 23.18 150.48 202.54 152.19 ;
   RECT 23.18 152.19 202.54 153.9 ;
   RECT 23.18 153.9 202.54 155.61 ;
   RECT 23.18 155.61 202.54 157.32 ;
   RECT 23.18 157.32 202.54 159.03 ;
   RECT 23.18 159.03 202.54 160.74 ;
   RECT 23.18 160.74 202.54 162.45 ;
   RECT 23.18 162.45 202.54 164.16 ;
   RECT 23.18 164.16 202.54 165.87 ;
   RECT 23.18 165.87 202.54 167.58 ;
   RECT 23.18 167.58 202.54 169.29 ;
   RECT 23.18 169.29 202.54 171.0 ;
   RECT 23.18 171.0 202.54 172.71 ;
   RECT 23.18 172.71 202.54 174.42 ;
   RECT 23.18 174.42 202.54 176.13 ;
   RECT 23.18 176.13 202.54 177.84 ;
   RECT 23.18 177.84 202.54 179.55 ;
   RECT 23.18 179.55 202.54 181.26 ;
   RECT 23.18 181.26 202.54 182.97 ;
   RECT 23.18 182.97 202.54 184.68 ;
   RECT 23.18 184.68 202.54 186.39 ;
   RECT 23.18 186.39 202.54 188.1 ;
   RECT 23.18 188.1 202.54 189.81 ;
   RECT 23.18 189.81 202.54 191.52 ;
   RECT 23.18 191.52 202.54 193.23 ;
   RECT 23.18 193.23 202.54 194.94 ;
   RECT 23.18 194.94 202.54 196.65 ;
   RECT 23.18 196.65 202.54 198.36 ;
   RECT 23.18 198.36 202.54 200.07 ;
   RECT 23.18 200.07 202.54 201.78 ;
   RECT 23.18 201.78 202.54 203.49 ;
   RECT 23.18 203.49 202.54 205.2 ;
   RECT 23.18 205.2 202.54 206.91 ;
   RECT 23.18 206.91 202.54 208.62 ;
   RECT 23.18 208.62 202.54 210.33 ;
   RECT 23.18 210.33 202.54 212.04 ;
   RECT 23.18 212.04 202.54 213.75 ;
   RECT 23.18 213.75 202.54 215.46 ;
   RECT 23.18 215.46 202.54 217.17 ;
   RECT 23.18 217.17 202.54 218.88 ;
   RECT 23.18 218.88 202.54 220.59 ;
   RECT 23.18 220.59 202.54 222.3 ;
   RECT 23.18 222.3 202.54 224.01 ;
   RECT 23.18 224.01 202.54 225.72 ;
   RECT 23.18 225.72 202.54 227.43 ;
   RECT 23.18 227.43 202.54 229.14 ;
   RECT 23.18 229.14 202.54 230.85 ;
   RECT 23.18 230.85 202.54 232.56 ;
   RECT 23.18 232.56 202.54 234.27 ;
   RECT 23.18 234.27 202.54 235.98 ;
   RECT 23.18 235.98 202.54 237.69 ;
   RECT 23.18 237.69 202.54 239.4 ;
   RECT 23.18 239.4 202.54 241.11 ;
   RECT 23.18 241.11 202.54 242.82 ;
   RECT 23.18 242.82 202.54 244.53 ;
   RECT 23.18 244.53 202.54 246.24 ;
   RECT 23.18 246.24 202.54 247.95 ;
   RECT 23.18 247.95 202.54 249.66 ;
   RECT 23.18 249.66 202.54 251.37 ;
   RECT 23.18 251.37 202.54 253.08 ;
   RECT 23.18 253.08 202.54 254.79 ;
   RECT 23.18 254.79 202.54 256.5 ;
   RECT 23.18 256.5 202.54 258.21 ;
   RECT 23.18 258.21 202.54 259.92 ;
   RECT 23.18 259.92 202.54 261.63 ;
   RECT 23.18 261.63 202.54 263.34 ;
   RECT 23.18 263.34 202.54 265.05 ;
   RECT 23.18 265.05 202.54 266.76 ;
   RECT 23.18 266.76 202.54 268.47 ;
   RECT 23.18 268.47 202.54 270.18 ;
   RECT 23.18 270.18 202.54 271.89 ;
   RECT 23.18 271.89 202.54 273.6 ;
   RECT 23.18 273.6 202.54 275.31 ;
   RECT 23.18 275.31 202.54 277.02 ;
   RECT 23.18 277.02 202.54 278.73 ;
   RECT 23.18 278.73 202.54 280.44 ;
   RECT 23.18 280.44 202.54 282.15 ;
   RECT 23.18 282.15 202.54 283.86 ;
   RECT 23.18 283.86 202.54 285.57 ;
   RECT 23.18 285.57 202.54 287.28 ;
   RECT 23.18 287.28 202.54 288.99 ;
   RECT 23.18 288.99 202.54 290.7 ;
   RECT 23.18 290.7 202.54 292.41 ;
   RECT 23.18 292.41 202.54 294.12 ;
   RECT 23.18 294.12 202.54 295.83 ;
   RECT 23.18 295.83 202.54 297.54 ;
   RECT 23.18 297.54 202.54 299.25 ;
   RECT 23.18 299.25 202.54 300.96 ;
   RECT 23.18 300.96 202.54 302.67 ;
   RECT 23.18 302.67 202.54 304.38 ;
   RECT 23.18 304.38 202.54 306.09 ;
   RECT 23.18 306.09 202.54 307.8 ;
   RECT 23.18 307.8 202.54 309.51 ;
   RECT 23.18 309.51 202.54 311.22 ;
   RECT 23.18 311.22 202.54 312.93 ;
   RECT 23.18 312.93 202.54 314.64 ;
   RECT 23.18 314.64 202.54 316.35 ;
   RECT 23.18 316.35 202.54 318.06 ;
   RECT 23.18 318.06 202.54 319.77 ;
   RECT 23.18 319.77 202.54 321.48 ;
   RECT 23.18 321.48 202.54 323.19 ;
   RECT 23.18 323.19 202.54 324.9 ;
   RECT 23.18 324.9 202.54 326.61 ;
   RECT 23.18 326.61 202.54 328.32 ;
   RECT 23.18 328.32 202.54 330.03 ;
   RECT 23.18 330.03 202.54 331.74 ;
   RECT 23.18 331.74 202.54 333.45 ;
   RECT 23.18 333.45 202.54 335.16 ;
   RECT 23.18 335.16 202.54 336.87 ;
   RECT 23.18 336.87 202.54 338.58 ;
   RECT 23.18 338.58 202.54 340.29 ;
   RECT 23.18 340.29 202.54 342.0 ;
   RECT 23.18 342.0 202.54 343.71 ;
   RECT 23.18 343.71 202.54 345.42 ;
   RECT 23.18 345.42 202.54 347.13 ;
   RECT 23.18 347.13 202.54 348.84 ;
   RECT 23.18 348.84 202.54 350.55 ;
   RECT 23.18 350.55 202.54 352.26 ;
   RECT 23.18 352.26 202.54 353.97 ;
   RECT 23.18 353.97 202.54 355.68 ;
   RECT 23.18 355.68 202.54 357.39 ;
   RECT 23.18 357.39 202.54 359.1 ;
   RECT 23.18 359.1 202.54 360.81 ;
   RECT 23.18 360.81 202.54 362.52 ;
   RECT 23.18 362.52 202.54 364.23 ;
   RECT 23.18 364.23 202.54 365.94 ;
   RECT 23.18 365.94 202.54 367.65 ;
   RECT 23.18 367.65 202.54 369.36 ;
   RECT 23.18 369.36 202.54 371.07 ;
   RECT 23.18 371.07 202.54 372.78 ;
   RECT 23.18 372.78 202.54 374.49 ;
   RECT 23.18 374.49 202.54 376.2 ;
   RECT 23.18 376.2 202.54 377.91 ;
   RECT 23.18 377.91 202.54 379.62 ;
   RECT 23.18 379.62 202.54 381.33 ;
   RECT 23.18 381.33 202.54 383.04 ;
   RECT 23.18 383.04 202.54 384.75 ;
   RECT 23.18 384.75 202.54 386.46 ;
   RECT 23.18 386.46 202.54 388.17 ;
   RECT 23.18 388.17 202.54 389.88 ;
   RECT 23.18 389.88 202.54 391.59 ;
   RECT 23.18 391.59 202.54 393.3 ;
   RECT 23.18 393.3 202.54 395.01 ;
   RECT 23.18 395.01 202.54 396.72 ;
   RECT 23.18 396.72 202.54 398.43 ;
   RECT 23.18 398.43 202.54 400.14 ;
   RECT 23.18 400.14 202.54 401.85 ;
   RECT 0.0 401.85 202.54 403.56 ;
   RECT 0.0 403.56 202.54 405.27 ;
   RECT 0.0 405.27 202.54 406.98 ;
   RECT 0.0 406.98 202.54 408.69 ;
   RECT 0.0 408.69 202.54 410.4 ;
   RECT 0.0 410.4 202.54 412.11 ;
   RECT 0.0 412.11 202.54 413.82 ;
   RECT 0.0 413.82 202.54 415.53 ;
   RECT 0.0 415.53 202.54 417.24 ;
   RECT 0.0 417.24 202.54 418.95 ;
   RECT 0.0 418.95 202.54 420.66 ;
   RECT 0.0 420.66 202.54 422.37 ;
   RECT 0.0 422.37 202.54 424.08 ;
   RECT 0.0 424.08 202.54 425.79 ;
   RECT 0.0 425.79 202.54 427.5 ;
   RECT 0.0 427.5 202.54 429.21 ;
   RECT 0.0 429.21 202.54 430.92 ;
   RECT 23.18 430.92 202.54 432.63 ;
   RECT 23.18 432.63 202.54 434.34 ;
   RECT 23.18 434.34 202.54 436.05 ;
   RECT 23.18 436.05 202.54 437.76 ;
   RECT 23.18 437.76 202.54 439.47 ;
   RECT 23.18 439.47 202.54 441.18 ;
   RECT 23.18 441.18 202.54 442.89 ;
   RECT 23.18 442.89 202.54 444.6 ;
   RECT 23.18 444.6 202.54 446.31 ;
   RECT 23.18 446.31 202.54 448.02 ;
   RECT 23.18 448.02 202.54 449.73 ;
   RECT 23.18 449.73 202.54 451.44 ;
   RECT 23.18 451.44 202.54 453.15 ;
   RECT 23.18 453.15 202.54 454.86 ;
   RECT 23.18 454.86 202.54 456.57 ;
   RECT 23.18 456.57 202.54 458.28 ;
   RECT 23.18 458.28 202.54 459.99 ;
   RECT 23.18 459.99 202.54 461.7 ;
   RECT 23.18 461.7 202.54 463.41 ;
   RECT 23.18 463.41 202.54 465.12 ;
   RECT 23.18 465.12 202.54 466.83 ;
   RECT 23.18 466.83 202.54 468.54 ;
   RECT 23.18 468.54 202.54 470.25 ;
   RECT 23.18 470.25 202.54 471.96 ;
   RECT 23.18 471.96 202.54 473.67 ;
   RECT 23.18 473.67 202.54 475.38 ;
   RECT 23.18 475.38 202.54 477.09 ;
   RECT 23.18 477.09 202.54 478.8 ;
   RECT 23.18 478.8 202.54 480.51 ;
   RECT 23.18 480.51 202.54 482.22 ;
   RECT 23.18 482.22 202.54 483.93 ;
   RECT 23.18 483.93 202.54 485.64 ;
   RECT 23.18 485.64 202.54 487.35 ;
   RECT 23.18 487.35 202.54 489.06 ;
   RECT 23.18 489.06 202.54 490.77 ;
   RECT 23.18 490.77 202.54 492.48 ;
   RECT 23.18 492.48 202.54 494.19 ;
   RECT 23.18 494.19 202.54 495.9 ;
   RECT 23.18 495.9 202.54 497.61 ;
   RECT 23.18 497.61 202.54 499.32 ;
   RECT 23.18 499.32 202.54 501.03 ;
   RECT 23.18 501.03 202.54 502.74 ;
   RECT 23.18 502.74 202.54 504.45 ;
   RECT 23.18 504.45 202.54 506.16 ;
   RECT 23.18 506.16 202.54 507.87 ;
   RECT 23.18 507.87 202.54 509.58 ;
   RECT 23.18 509.58 202.54 511.29 ;
   RECT 23.18 511.29 202.54 513.0 ;
   RECT 23.18 513.0 202.54 514.71 ;
   RECT 23.18 514.71 202.54 516.42 ;
   RECT 23.18 516.42 202.54 518.13 ;
   RECT 23.18 518.13 202.54 519.84 ;
   RECT 23.18 519.84 202.54 521.55 ;
   RECT 23.18 521.55 202.54 523.26 ;
   RECT 23.18 523.26 202.54 524.97 ;
   RECT 23.18 524.97 202.54 526.68 ;
   RECT 23.18 526.68 202.54 528.39 ;
   RECT 23.18 528.39 202.54 530.1 ;
   RECT 23.18 530.1 202.54 531.81 ;
   RECT 23.18 531.81 202.54 533.52 ;
   RECT 23.18 533.52 202.54 535.23 ;
   RECT 23.18 535.23 202.54 536.94 ;
   RECT 23.18 536.94 202.54 538.65 ;
   RECT 23.18 538.65 202.54 540.36 ;
   RECT 23.18 540.36 202.54 542.07 ;
   RECT 23.18 542.07 202.54 543.78 ;
   RECT 23.18 543.78 202.54 545.49 ;
   RECT 23.18 545.49 202.54 547.2 ;
   RECT 23.18 547.2 202.54 548.91 ;
   RECT 23.18 548.91 202.54 550.62 ;
   RECT 23.18 550.62 202.54 552.33 ;
   RECT 23.18 552.33 202.54 554.04 ;
   RECT 23.18 554.04 202.54 555.75 ;
   RECT 23.18 555.75 202.54 557.46 ;
   RECT 23.18 557.46 202.54 559.17 ;
   RECT 23.18 559.17 202.54 560.88 ;
   RECT 23.18 560.88 202.54 562.59 ;
   RECT 23.18 562.59 202.54 564.3 ;
   RECT 23.18 564.3 202.54 566.01 ;
   RECT 23.18 566.01 202.54 567.72 ;
   RECT 23.18 567.72 202.54 569.43 ;
   RECT 23.18 569.43 202.54 571.14 ;
   RECT 23.18 571.14 202.54 572.85 ;
   RECT 23.18 572.85 202.54 574.56 ;
   RECT 23.18 574.56 202.54 576.27 ;
   RECT 23.18 576.27 202.54 577.98 ;
   RECT 23.18 577.98 202.54 579.69 ;
   RECT 23.18 579.69 202.54 581.4 ;
   RECT 23.18 581.4 202.54 583.11 ;
   RECT 23.18 583.11 202.54 584.82 ;
   RECT 23.18 584.82 202.54 586.53 ;
   RECT 23.18 586.53 202.54 588.24 ;
   RECT 23.18 588.24 202.54 589.95 ;
   RECT 23.18 589.95 202.54 591.66 ;
   RECT 23.18 591.66 202.54 593.37 ;
   RECT 23.18 593.37 202.54 595.08 ;
   RECT 23.18 595.08 202.54 596.79 ;
   RECT 23.18 596.79 202.54 598.5 ;
   RECT 23.18 598.5 202.54 600.21 ;
   RECT 23.18 600.21 202.54 601.92 ;
   RECT 23.18 601.92 202.54 603.63 ;
   RECT 23.18 603.63 202.54 605.34 ;
   RECT 23.18 605.34 202.54 607.05 ;
   RECT 23.18 607.05 202.54 608.76 ;
   RECT 23.18 608.76 202.54 610.47 ;
   RECT 23.18 610.47 202.54 612.18 ;
   RECT 23.18 612.18 202.54 613.89 ;
   RECT 23.18 613.89 202.54 615.6 ;
   RECT 23.18 615.6 202.54 617.31 ;
   RECT 23.18 617.31 202.54 619.02 ;
   RECT 23.18 619.02 202.54 620.73 ;
   RECT 23.18 620.73 202.54 622.44 ;
   RECT 23.18 622.44 202.54 624.15 ;
   RECT 23.18 624.15 202.54 625.86 ;
   RECT 23.18 625.86 202.54 627.57 ;
   RECT 23.18 627.57 202.54 629.28 ;
   RECT 23.18 629.28 202.54 630.99 ;
   RECT 23.18 630.99 202.54 632.7 ;
   RECT 23.18 632.7 202.54 634.41 ;
   RECT 23.18 634.41 202.54 636.12 ;
   RECT 23.18 636.12 202.54 637.83 ;
   RECT 23.18 637.83 202.54 639.54 ;
   RECT 23.18 639.54 202.54 641.25 ;
   RECT 23.18 641.25 202.54 642.96 ;
   RECT 23.18 642.96 202.54 644.67 ;
   RECT 23.18 644.67 202.54 646.38 ;
   RECT 23.18 646.38 202.54 648.09 ;
   RECT 23.18 648.09 202.54 649.8 ;
   RECT 23.18 649.8 202.54 651.51 ;
   RECT 23.18 651.51 202.54 653.22 ;
   RECT 23.18 653.22 202.54 654.93 ;
   RECT 23.18 654.93 202.54 656.64 ;
   RECT 23.18 656.64 202.54 658.35 ;
   RECT 23.18 658.35 202.54 660.06 ;
   RECT 23.18 660.06 202.54 661.77 ;
   RECT 23.18 661.77 202.54 663.48 ;
   RECT 23.18 663.48 202.54 665.19 ;
   RECT 23.18 665.19 202.54 666.9 ;
   RECT 23.18 666.9 202.54 668.61 ;
   RECT 23.18 668.61 202.54 670.32 ;
   RECT 23.18 670.32 202.54 672.03 ;
   RECT 23.18 672.03 202.54 673.74 ;
   RECT 23.18 673.74 202.54 675.45 ;
   RECT 23.18 675.45 202.54 677.16 ;
   RECT 23.18 677.16 202.54 678.87 ;
   RECT 23.18 678.87 202.54 680.58 ;
   RECT 23.18 680.58 202.54 682.29 ;
   RECT 23.18 682.29 202.54 684.0 ;
   RECT 23.18 684.0 202.54 685.71 ;
   RECT 23.18 685.71 202.54 687.42 ;
   RECT 23.18 687.42 202.54 689.13 ;
   RECT 23.18 689.13 202.54 690.84 ;
   RECT 23.18 690.84 202.54 692.55 ;
   RECT 23.18 692.55 202.54 694.26 ;
   RECT 23.18 694.26 202.54 695.97 ;
   RECT 23.18 695.97 202.54 697.68 ;
   RECT 23.18 697.68 202.54 699.39 ;
   RECT 23.18 699.39 202.54 701.1 ;
   RECT 23.18 701.1 202.54 702.81 ;
   RECT 23.18 702.81 202.54 704.52 ;
   RECT 23.18 704.52 202.54 706.23 ;
   RECT 23.18 706.23 202.54 707.94 ;
   RECT 23.18 707.94 202.54 709.65 ;
   RECT 23.18 709.65 202.54 711.36 ;
   RECT 23.18 711.36 202.54 713.07 ;
   RECT 23.18 713.07 202.54 714.78 ;
   RECT 23.18 714.78 202.54 716.49 ;
   RECT 23.18 716.49 202.54 718.2 ;
   RECT 23.18 718.2 202.54 719.91 ;
   RECT 23.18 719.91 202.54 721.62 ;
   RECT 23.18 721.62 202.54 723.33 ;
   RECT 23.18 723.33 202.54 725.04 ;
   RECT 23.18 725.04 202.54 726.75 ;
   RECT 23.18 726.75 202.54 728.46 ;
   RECT 23.18 728.46 202.54 730.17 ;
   RECT 23.18 730.17 202.54 731.88 ;
   RECT 23.18 731.88 202.54 733.59 ;
   RECT 23.18 733.59 202.54 735.3 ;
   RECT 23.18 735.3 202.54 737.01 ;
   RECT 23.18 737.01 202.54 738.72 ;
   RECT 23.18 738.72 202.54 740.43 ;
   RECT 23.18 740.43 202.54 742.14 ;
   RECT 23.18 742.14 202.54 743.85 ;
   RECT 23.18 743.85 202.54 745.56 ;
   RECT 23.18 745.56 202.54 747.27 ;
   RECT 23.18 747.27 202.54 748.98 ;
   RECT 23.18 748.98 202.54 750.69 ;
   RECT 23.18 750.69 202.54 752.4 ;
   RECT 23.18 752.4 202.54 754.11 ;
   RECT 23.18 754.11 202.54 755.82 ;
   RECT 23.18 755.82 202.54 757.53 ;
   RECT 23.18 757.53 202.54 759.24 ;
   RECT 23.18 759.24 202.54 760.95 ;
   RECT 23.18 760.95 202.54 762.66 ;
   RECT 23.18 762.66 202.54 764.37 ;
   RECT 23.18 764.37 202.54 766.08 ;
   RECT 23.18 766.08 202.54 767.79 ;
   RECT 23.18 767.79 202.54 769.5 ;
   RECT 23.18 769.5 202.54 771.21 ;
   RECT 23.18 771.21 202.54 772.92 ;
   RECT 23.18 772.92 202.54 774.63 ;
   RECT 23.18 774.63 202.54 776.34 ;
   RECT 23.18 776.34 202.54 778.05 ;
   RECT 23.18 778.05 202.54 779.76 ;
   RECT 23.18 779.76 202.54 781.47 ;
   RECT 23.18 781.47 202.54 783.18 ;
   RECT 23.18 783.18 202.54 784.89 ;
   RECT 23.18 784.89 202.54 786.6 ;
   RECT 23.18 786.6 202.54 788.31 ;
   RECT 23.18 788.31 202.54 790.02 ;
   RECT 23.18 790.02 202.54 791.73 ;
   RECT 23.18 791.73 202.54 793.44 ;
   RECT 23.18 793.44 202.54 795.15 ;
   RECT 23.18 795.15 202.54 796.86 ;
   RECT 23.18 796.86 202.54 798.57 ;
   RECT 23.18 798.57 202.54 800.28 ;
   RECT 23.18 800.28 202.54 801.99 ;
   RECT 23.18 801.99 202.54 803.7 ;
   RECT 23.18 803.7 202.54 805.41 ;
   RECT 23.18 805.41 202.54 807.12 ;
   RECT 23.18 807.12 202.54 808.83 ;
   RECT 23.18 808.83 202.54 810.54 ;
   RECT 23.18 810.54 202.54 812.25 ;
   RECT 23.18 812.25 202.54 813.96 ;
   RECT 23.18 813.96 202.54 815.67 ;
   RECT 23.18 815.67 202.54 817.38 ;
   RECT 23.18 817.38 202.54 819.09 ;
   RECT 23.18 819.09 202.54 820.8 ;
   RECT 23.18 820.8 202.54 822.51 ;
   RECT 23.18 822.51 202.54 824.22 ;
   RECT 23.18 824.22 202.54 825.93 ;
   RECT 23.18 825.93 202.54 827.64 ;
   RECT 23.18 827.64 202.54 829.35 ;
   RECT 23.18 829.35 202.54 831.06 ;
   RECT 23.18 831.06 202.54 832.77 ;
   RECT 23.18 832.77 202.54 834.48 ;
   RECT 23.18 834.48 202.54 836.19 ;
   RECT 23.18 836.19 202.54 837.9 ;
   RECT 23.18 837.9 202.54 839.61 ;
   RECT 23.18 839.61 202.54 841.32 ;
  LAYER metal2 ;
   RECT 23.18 0.0 202.54 1.71 ;
   RECT 23.18 1.71 202.54 3.42 ;
   RECT 23.18 3.42 202.54 5.13 ;
   RECT 23.18 5.13 202.54 6.84 ;
   RECT 23.18 6.84 202.54 8.55 ;
   RECT 23.18 8.55 202.54 10.26 ;
   RECT 23.18 10.26 202.54 11.97 ;
   RECT 23.18 11.97 202.54 13.68 ;
   RECT 23.18 13.68 202.54 15.39 ;
   RECT 23.18 15.39 202.54 17.1 ;
   RECT 23.18 17.1 202.54 18.81 ;
   RECT 23.18 18.81 202.54 20.52 ;
   RECT 23.18 20.52 202.54 22.23 ;
   RECT 23.18 22.23 202.54 23.94 ;
   RECT 23.18 23.94 202.54 25.65 ;
   RECT 23.18 25.65 202.54 27.36 ;
   RECT 23.18 27.36 202.54 29.07 ;
   RECT 23.18 29.07 202.54 30.78 ;
   RECT 23.18 30.78 202.54 32.49 ;
   RECT 23.18 32.49 202.54 34.2 ;
   RECT 23.18 34.2 202.54 35.91 ;
   RECT 23.18 35.91 202.54 37.62 ;
   RECT 23.18 37.62 202.54 39.33 ;
   RECT 23.18 39.33 202.54 41.04 ;
   RECT 23.18 41.04 202.54 42.75 ;
   RECT 23.18 42.75 202.54 44.46 ;
   RECT 23.18 44.46 202.54 46.17 ;
   RECT 23.18 46.17 202.54 47.88 ;
   RECT 23.18 47.88 202.54 49.59 ;
   RECT 23.18 49.59 202.54 51.3 ;
   RECT 23.18 51.3 202.54 53.01 ;
   RECT 23.18 53.01 202.54 54.72 ;
   RECT 23.18 54.72 202.54 56.43 ;
   RECT 23.18 56.43 202.54 58.14 ;
   RECT 23.18 58.14 202.54 59.85 ;
   RECT 23.18 59.85 202.54 61.56 ;
   RECT 23.18 61.56 202.54 63.27 ;
   RECT 23.18 63.27 202.54 64.98 ;
   RECT 23.18 64.98 202.54 66.69 ;
   RECT 23.18 66.69 202.54 68.4 ;
   RECT 23.18 68.4 202.54 70.11 ;
   RECT 23.18 70.11 202.54 71.82 ;
   RECT 23.18 71.82 202.54 73.53 ;
   RECT 23.18 73.53 202.54 75.24 ;
   RECT 23.18 75.24 202.54 76.95 ;
   RECT 23.18 76.95 202.54 78.66 ;
   RECT 23.18 78.66 202.54 80.37 ;
   RECT 23.18 80.37 202.54 82.08 ;
   RECT 23.18 82.08 202.54 83.79 ;
   RECT 23.18 83.79 202.54 85.5 ;
   RECT 23.18 85.5 202.54 87.21 ;
   RECT 23.18 87.21 202.54 88.92 ;
   RECT 23.18 88.92 202.54 90.63 ;
   RECT 23.18 90.63 202.54 92.34 ;
   RECT 23.18 92.34 202.54 94.05 ;
   RECT 23.18 94.05 202.54 95.76 ;
   RECT 23.18 95.76 202.54 97.47 ;
   RECT 23.18 97.47 202.54 99.18 ;
   RECT 23.18 99.18 202.54 100.89 ;
   RECT 23.18 100.89 202.54 102.6 ;
   RECT 23.18 102.6 202.54 104.31 ;
   RECT 23.18 104.31 202.54 106.02 ;
   RECT 23.18 106.02 202.54 107.73 ;
   RECT 23.18 107.73 202.54 109.44 ;
   RECT 23.18 109.44 202.54 111.15 ;
   RECT 23.18 111.15 202.54 112.86 ;
   RECT 23.18 112.86 202.54 114.57 ;
   RECT 23.18 114.57 202.54 116.28 ;
   RECT 23.18 116.28 202.54 117.99 ;
   RECT 23.18 117.99 202.54 119.7 ;
   RECT 23.18 119.7 202.54 121.41 ;
   RECT 23.18 121.41 202.54 123.12 ;
   RECT 23.18 123.12 202.54 124.83 ;
   RECT 23.18 124.83 202.54 126.54 ;
   RECT 23.18 126.54 202.54 128.25 ;
   RECT 23.18 128.25 202.54 129.96 ;
   RECT 23.18 129.96 202.54 131.67 ;
   RECT 23.18 131.67 202.54 133.38 ;
   RECT 23.18 133.38 202.54 135.09 ;
   RECT 23.18 135.09 202.54 136.8 ;
   RECT 23.18 136.8 202.54 138.51 ;
   RECT 23.18 138.51 202.54 140.22 ;
   RECT 23.18 140.22 202.54 141.93 ;
   RECT 23.18 141.93 202.54 143.64 ;
   RECT 23.18 143.64 202.54 145.35 ;
   RECT 23.18 145.35 202.54 147.06 ;
   RECT 23.18 147.06 202.54 148.77 ;
   RECT 23.18 148.77 202.54 150.48 ;
   RECT 23.18 150.48 202.54 152.19 ;
   RECT 23.18 152.19 202.54 153.9 ;
   RECT 23.18 153.9 202.54 155.61 ;
   RECT 23.18 155.61 202.54 157.32 ;
   RECT 23.18 157.32 202.54 159.03 ;
   RECT 23.18 159.03 202.54 160.74 ;
   RECT 23.18 160.74 202.54 162.45 ;
   RECT 23.18 162.45 202.54 164.16 ;
   RECT 23.18 164.16 202.54 165.87 ;
   RECT 23.18 165.87 202.54 167.58 ;
   RECT 23.18 167.58 202.54 169.29 ;
   RECT 23.18 169.29 202.54 171.0 ;
   RECT 23.18 171.0 202.54 172.71 ;
   RECT 23.18 172.71 202.54 174.42 ;
   RECT 23.18 174.42 202.54 176.13 ;
   RECT 23.18 176.13 202.54 177.84 ;
   RECT 23.18 177.84 202.54 179.55 ;
   RECT 23.18 179.55 202.54 181.26 ;
   RECT 23.18 181.26 202.54 182.97 ;
   RECT 23.18 182.97 202.54 184.68 ;
   RECT 23.18 184.68 202.54 186.39 ;
   RECT 23.18 186.39 202.54 188.1 ;
   RECT 23.18 188.1 202.54 189.81 ;
   RECT 23.18 189.81 202.54 191.52 ;
   RECT 23.18 191.52 202.54 193.23 ;
   RECT 23.18 193.23 202.54 194.94 ;
   RECT 23.18 194.94 202.54 196.65 ;
   RECT 23.18 196.65 202.54 198.36 ;
   RECT 23.18 198.36 202.54 200.07 ;
   RECT 23.18 200.07 202.54 201.78 ;
   RECT 23.18 201.78 202.54 203.49 ;
   RECT 23.18 203.49 202.54 205.2 ;
   RECT 23.18 205.2 202.54 206.91 ;
   RECT 23.18 206.91 202.54 208.62 ;
   RECT 23.18 208.62 202.54 210.33 ;
   RECT 23.18 210.33 202.54 212.04 ;
   RECT 23.18 212.04 202.54 213.75 ;
   RECT 23.18 213.75 202.54 215.46 ;
   RECT 23.18 215.46 202.54 217.17 ;
   RECT 23.18 217.17 202.54 218.88 ;
   RECT 23.18 218.88 202.54 220.59 ;
   RECT 23.18 220.59 202.54 222.3 ;
   RECT 23.18 222.3 202.54 224.01 ;
   RECT 23.18 224.01 202.54 225.72 ;
   RECT 23.18 225.72 202.54 227.43 ;
   RECT 23.18 227.43 202.54 229.14 ;
   RECT 23.18 229.14 202.54 230.85 ;
   RECT 23.18 230.85 202.54 232.56 ;
   RECT 23.18 232.56 202.54 234.27 ;
   RECT 23.18 234.27 202.54 235.98 ;
   RECT 23.18 235.98 202.54 237.69 ;
   RECT 23.18 237.69 202.54 239.4 ;
   RECT 23.18 239.4 202.54 241.11 ;
   RECT 23.18 241.11 202.54 242.82 ;
   RECT 23.18 242.82 202.54 244.53 ;
   RECT 23.18 244.53 202.54 246.24 ;
   RECT 23.18 246.24 202.54 247.95 ;
   RECT 23.18 247.95 202.54 249.66 ;
   RECT 23.18 249.66 202.54 251.37 ;
   RECT 23.18 251.37 202.54 253.08 ;
   RECT 23.18 253.08 202.54 254.79 ;
   RECT 23.18 254.79 202.54 256.5 ;
   RECT 23.18 256.5 202.54 258.21 ;
   RECT 23.18 258.21 202.54 259.92 ;
   RECT 23.18 259.92 202.54 261.63 ;
   RECT 23.18 261.63 202.54 263.34 ;
   RECT 23.18 263.34 202.54 265.05 ;
   RECT 23.18 265.05 202.54 266.76 ;
   RECT 23.18 266.76 202.54 268.47 ;
   RECT 23.18 268.47 202.54 270.18 ;
   RECT 23.18 270.18 202.54 271.89 ;
   RECT 23.18 271.89 202.54 273.6 ;
   RECT 23.18 273.6 202.54 275.31 ;
   RECT 23.18 275.31 202.54 277.02 ;
   RECT 23.18 277.02 202.54 278.73 ;
   RECT 23.18 278.73 202.54 280.44 ;
   RECT 23.18 280.44 202.54 282.15 ;
   RECT 23.18 282.15 202.54 283.86 ;
   RECT 23.18 283.86 202.54 285.57 ;
   RECT 23.18 285.57 202.54 287.28 ;
   RECT 23.18 287.28 202.54 288.99 ;
   RECT 23.18 288.99 202.54 290.7 ;
   RECT 23.18 290.7 202.54 292.41 ;
   RECT 23.18 292.41 202.54 294.12 ;
   RECT 23.18 294.12 202.54 295.83 ;
   RECT 23.18 295.83 202.54 297.54 ;
   RECT 23.18 297.54 202.54 299.25 ;
   RECT 23.18 299.25 202.54 300.96 ;
   RECT 23.18 300.96 202.54 302.67 ;
   RECT 23.18 302.67 202.54 304.38 ;
   RECT 23.18 304.38 202.54 306.09 ;
   RECT 23.18 306.09 202.54 307.8 ;
   RECT 23.18 307.8 202.54 309.51 ;
   RECT 23.18 309.51 202.54 311.22 ;
   RECT 23.18 311.22 202.54 312.93 ;
   RECT 23.18 312.93 202.54 314.64 ;
   RECT 23.18 314.64 202.54 316.35 ;
   RECT 23.18 316.35 202.54 318.06 ;
   RECT 23.18 318.06 202.54 319.77 ;
   RECT 23.18 319.77 202.54 321.48 ;
   RECT 23.18 321.48 202.54 323.19 ;
   RECT 23.18 323.19 202.54 324.9 ;
   RECT 23.18 324.9 202.54 326.61 ;
   RECT 23.18 326.61 202.54 328.32 ;
   RECT 23.18 328.32 202.54 330.03 ;
   RECT 23.18 330.03 202.54 331.74 ;
   RECT 23.18 331.74 202.54 333.45 ;
   RECT 23.18 333.45 202.54 335.16 ;
   RECT 23.18 335.16 202.54 336.87 ;
   RECT 23.18 336.87 202.54 338.58 ;
   RECT 23.18 338.58 202.54 340.29 ;
   RECT 23.18 340.29 202.54 342.0 ;
   RECT 23.18 342.0 202.54 343.71 ;
   RECT 23.18 343.71 202.54 345.42 ;
   RECT 23.18 345.42 202.54 347.13 ;
   RECT 23.18 347.13 202.54 348.84 ;
   RECT 23.18 348.84 202.54 350.55 ;
   RECT 23.18 350.55 202.54 352.26 ;
   RECT 23.18 352.26 202.54 353.97 ;
   RECT 23.18 353.97 202.54 355.68 ;
   RECT 23.18 355.68 202.54 357.39 ;
   RECT 23.18 357.39 202.54 359.1 ;
   RECT 23.18 359.1 202.54 360.81 ;
   RECT 23.18 360.81 202.54 362.52 ;
   RECT 23.18 362.52 202.54 364.23 ;
   RECT 23.18 364.23 202.54 365.94 ;
   RECT 23.18 365.94 202.54 367.65 ;
   RECT 23.18 367.65 202.54 369.36 ;
   RECT 23.18 369.36 202.54 371.07 ;
   RECT 23.18 371.07 202.54 372.78 ;
   RECT 23.18 372.78 202.54 374.49 ;
   RECT 23.18 374.49 202.54 376.2 ;
   RECT 23.18 376.2 202.54 377.91 ;
   RECT 23.18 377.91 202.54 379.62 ;
   RECT 23.18 379.62 202.54 381.33 ;
   RECT 23.18 381.33 202.54 383.04 ;
   RECT 23.18 383.04 202.54 384.75 ;
   RECT 23.18 384.75 202.54 386.46 ;
   RECT 23.18 386.46 202.54 388.17 ;
   RECT 23.18 388.17 202.54 389.88 ;
   RECT 23.18 389.88 202.54 391.59 ;
   RECT 23.18 391.59 202.54 393.3 ;
   RECT 23.18 393.3 202.54 395.01 ;
   RECT 23.18 395.01 202.54 396.72 ;
   RECT 23.18 396.72 202.54 398.43 ;
   RECT 23.18 398.43 202.54 400.14 ;
   RECT 23.18 400.14 202.54 401.85 ;
   RECT 0.0 401.85 202.54 403.56 ;
   RECT 0.0 403.56 202.54 405.27 ;
   RECT 0.0 405.27 202.54 406.98 ;
   RECT 0.0 406.98 202.54 408.69 ;
   RECT 0.0 408.69 202.54 410.4 ;
   RECT 0.0 410.4 202.54 412.11 ;
   RECT 0.0 412.11 202.54 413.82 ;
   RECT 0.0 413.82 202.54 415.53 ;
   RECT 0.0 415.53 202.54 417.24 ;
   RECT 0.0 417.24 202.54 418.95 ;
   RECT 0.0 418.95 202.54 420.66 ;
   RECT 0.0 420.66 202.54 422.37 ;
   RECT 0.0 422.37 202.54 424.08 ;
   RECT 0.0 424.08 202.54 425.79 ;
   RECT 0.0 425.79 202.54 427.5 ;
   RECT 0.0 427.5 202.54 429.21 ;
   RECT 0.0 429.21 202.54 430.92 ;
   RECT 23.18 430.92 202.54 432.63 ;
   RECT 23.18 432.63 202.54 434.34 ;
   RECT 23.18 434.34 202.54 436.05 ;
   RECT 23.18 436.05 202.54 437.76 ;
   RECT 23.18 437.76 202.54 439.47 ;
   RECT 23.18 439.47 202.54 441.18 ;
   RECT 23.18 441.18 202.54 442.89 ;
   RECT 23.18 442.89 202.54 444.6 ;
   RECT 23.18 444.6 202.54 446.31 ;
   RECT 23.18 446.31 202.54 448.02 ;
   RECT 23.18 448.02 202.54 449.73 ;
   RECT 23.18 449.73 202.54 451.44 ;
   RECT 23.18 451.44 202.54 453.15 ;
   RECT 23.18 453.15 202.54 454.86 ;
   RECT 23.18 454.86 202.54 456.57 ;
   RECT 23.18 456.57 202.54 458.28 ;
   RECT 23.18 458.28 202.54 459.99 ;
   RECT 23.18 459.99 202.54 461.7 ;
   RECT 23.18 461.7 202.54 463.41 ;
   RECT 23.18 463.41 202.54 465.12 ;
   RECT 23.18 465.12 202.54 466.83 ;
   RECT 23.18 466.83 202.54 468.54 ;
   RECT 23.18 468.54 202.54 470.25 ;
   RECT 23.18 470.25 202.54 471.96 ;
   RECT 23.18 471.96 202.54 473.67 ;
   RECT 23.18 473.67 202.54 475.38 ;
   RECT 23.18 475.38 202.54 477.09 ;
   RECT 23.18 477.09 202.54 478.8 ;
   RECT 23.18 478.8 202.54 480.51 ;
   RECT 23.18 480.51 202.54 482.22 ;
   RECT 23.18 482.22 202.54 483.93 ;
   RECT 23.18 483.93 202.54 485.64 ;
   RECT 23.18 485.64 202.54 487.35 ;
   RECT 23.18 487.35 202.54 489.06 ;
   RECT 23.18 489.06 202.54 490.77 ;
   RECT 23.18 490.77 202.54 492.48 ;
   RECT 23.18 492.48 202.54 494.19 ;
   RECT 23.18 494.19 202.54 495.9 ;
   RECT 23.18 495.9 202.54 497.61 ;
   RECT 23.18 497.61 202.54 499.32 ;
   RECT 23.18 499.32 202.54 501.03 ;
   RECT 23.18 501.03 202.54 502.74 ;
   RECT 23.18 502.74 202.54 504.45 ;
   RECT 23.18 504.45 202.54 506.16 ;
   RECT 23.18 506.16 202.54 507.87 ;
   RECT 23.18 507.87 202.54 509.58 ;
   RECT 23.18 509.58 202.54 511.29 ;
   RECT 23.18 511.29 202.54 513.0 ;
   RECT 23.18 513.0 202.54 514.71 ;
   RECT 23.18 514.71 202.54 516.42 ;
   RECT 23.18 516.42 202.54 518.13 ;
   RECT 23.18 518.13 202.54 519.84 ;
   RECT 23.18 519.84 202.54 521.55 ;
   RECT 23.18 521.55 202.54 523.26 ;
   RECT 23.18 523.26 202.54 524.97 ;
   RECT 23.18 524.97 202.54 526.68 ;
   RECT 23.18 526.68 202.54 528.39 ;
   RECT 23.18 528.39 202.54 530.1 ;
   RECT 23.18 530.1 202.54 531.81 ;
   RECT 23.18 531.81 202.54 533.52 ;
   RECT 23.18 533.52 202.54 535.23 ;
   RECT 23.18 535.23 202.54 536.94 ;
   RECT 23.18 536.94 202.54 538.65 ;
   RECT 23.18 538.65 202.54 540.36 ;
   RECT 23.18 540.36 202.54 542.07 ;
   RECT 23.18 542.07 202.54 543.78 ;
   RECT 23.18 543.78 202.54 545.49 ;
   RECT 23.18 545.49 202.54 547.2 ;
   RECT 23.18 547.2 202.54 548.91 ;
   RECT 23.18 548.91 202.54 550.62 ;
   RECT 23.18 550.62 202.54 552.33 ;
   RECT 23.18 552.33 202.54 554.04 ;
   RECT 23.18 554.04 202.54 555.75 ;
   RECT 23.18 555.75 202.54 557.46 ;
   RECT 23.18 557.46 202.54 559.17 ;
   RECT 23.18 559.17 202.54 560.88 ;
   RECT 23.18 560.88 202.54 562.59 ;
   RECT 23.18 562.59 202.54 564.3 ;
   RECT 23.18 564.3 202.54 566.01 ;
   RECT 23.18 566.01 202.54 567.72 ;
   RECT 23.18 567.72 202.54 569.43 ;
   RECT 23.18 569.43 202.54 571.14 ;
   RECT 23.18 571.14 202.54 572.85 ;
   RECT 23.18 572.85 202.54 574.56 ;
   RECT 23.18 574.56 202.54 576.27 ;
   RECT 23.18 576.27 202.54 577.98 ;
   RECT 23.18 577.98 202.54 579.69 ;
   RECT 23.18 579.69 202.54 581.4 ;
   RECT 23.18 581.4 202.54 583.11 ;
   RECT 23.18 583.11 202.54 584.82 ;
   RECT 23.18 584.82 202.54 586.53 ;
   RECT 23.18 586.53 202.54 588.24 ;
   RECT 23.18 588.24 202.54 589.95 ;
   RECT 23.18 589.95 202.54 591.66 ;
   RECT 23.18 591.66 202.54 593.37 ;
   RECT 23.18 593.37 202.54 595.08 ;
   RECT 23.18 595.08 202.54 596.79 ;
   RECT 23.18 596.79 202.54 598.5 ;
   RECT 23.18 598.5 202.54 600.21 ;
   RECT 23.18 600.21 202.54 601.92 ;
   RECT 23.18 601.92 202.54 603.63 ;
   RECT 23.18 603.63 202.54 605.34 ;
   RECT 23.18 605.34 202.54 607.05 ;
   RECT 23.18 607.05 202.54 608.76 ;
   RECT 23.18 608.76 202.54 610.47 ;
   RECT 23.18 610.47 202.54 612.18 ;
   RECT 23.18 612.18 202.54 613.89 ;
   RECT 23.18 613.89 202.54 615.6 ;
   RECT 23.18 615.6 202.54 617.31 ;
   RECT 23.18 617.31 202.54 619.02 ;
   RECT 23.18 619.02 202.54 620.73 ;
   RECT 23.18 620.73 202.54 622.44 ;
   RECT 23.18 622.44 202.54 624.15 ;
   RECT 23.18 624.15 202.54 625.86 ;
   RECT 23.18 625.86 202.54 627.57 ;
   RECT 23.18 627.57 202.54 629.28 ;
   RECT 23.18 629.28 202.54 630.99 ;
   RECT 23.18 630.99 202.54 632.7 ;
   RECT 23.18 632.7 202.54 634.41 ;
   RECT 23.18 634.41 202.54 636.12 ;
   RECT 23.18 636.12 202.54 637.83 ;
   RECT 23.18 637.83 202.54 639.54 ;
   RECT 23.18 639.54 202.54 641.25 ;
   RECT 23.18 641.25 202.54 642.96 ;
   RECT 23.18 642.96 202.54 644.67 ;
   RECT 23.18 644.67 202.54 646.38 ;
   RECT 23.18 646.38 202.54 648.09 ;
   RECT 23.18 648.09 202.54 649.8 ;
   RECT 23.18 649.8 202.54 651.51 ;
   RECT 23.18 651.51 202.54 653.22 ;
   RECT 23.18 653.22 202.54 654.93 ;
   RECT 23.18 654.93 202.54 656.64 ;
   RECT 23.18 656.64 202.54 658.35 ;
   RECT 23.18 658.35 202.54 660.06 ;
   RECT 23.18 660.06 202.54 661.77 ;
   RECT 23.18 661.77 202.54 663.48 ;
   RECT 23.18 663.48 202.54 665.19 ;
   RECT 23.18 665.19 202.54 666.9 ;
   RECT 23.18 666.9 202.54 668.61 ;
   RECT 23.18 668.61 202.54 670.32 ;
   RECT 23.18 670.32 202.54 672.03 ;
   RECT 23.18 672.03 202.54 673.74 ;
   RECT 23.18 673.74 202.54 675.45 ;
   RECT 23.18 675.45 202.54 677.16 ;
   RECT 23.18 677.16 202.54 678.87 ;
   RECT 23.18 678.87 202.54 680.58 ;
   RECT 23.18 680.58 202.54 682.29 ;
   RECT 23.18 682.29 202.54 684.0 ;
   RECT 23.18 684.0 202.54 685.71 ;
   RECT 23.18 685.71 202.54 687.42 ;
   RECT 23.18 687.42 202.54 689.13 ;
   RECT 23.18 689.13 202.54 690.84 ;
   RECT 23.18 690.84 202.54 692.55 ;
   RECT 23.18 692.55 202.54 694.26 ;
   RECT 23.18 694.26 202.54 695.97 ;
   RECT 23.18 695.97 202.54 697.68 ;
   RECT 23.18 697.68 202.54 699.39 ;
   RECT 23.18 699.39 202.54 701.1 ;
   RECT 23.18 701.1 202.54 702.81 ;
   RECT 23.18 702.81 202.54 704.52 ;
   RECT 23.18 704.52 202.54 706.23 ;
   RECT 23.18 706.23 202.54 707.94 ;
   RECT 23.18 707.94 202.54 709.65 ;
   RECT 23.18 709.65 202.54 711.36 ;
   RECT 23.18 711.36 202.54 713.07 ;
   RECT 23.18 713.07 202.54 714.78 ;
   RECT 23.18 714.78 202.54 716.49 ;
   RECT 23.18 716.49 202.54 718.2 ;
   RECT 23.18 718.2 202.54 719.91 ;
   RECT 23.18 719.91 202.54 721.62 ;
   RECT 23.18 721.62 202.54 723.33 ;
   RECT 23.18 723.33 202.54 725.04 ;
   RECT 23.18 725.04 202.54 726.75 ;
   RECT 23.18 726.75 202.54 728.46 ;
   RECT 23.18 728.46 202.54 730.17 ;
   RECT 23.18 730.17 202.54 731.88 ;
   RECT 23.18 731.88 202.54 733.59 ;
   RECT 23.18 733.59 202.54 735.3 ;
   RECT 23.18 735.3 202.54 737.01 ;
   RECT 23.18 737.01 202.54 738.72 ;
   RECT 23.18 738.72 202.54 740.43 ;
   RECT 23.18 740.43 202.54 742.14 ;
   RECT 23.18 742.14 202.54 743.85 ;
   RECT 23.18 743.85 202.54 745.56 ;
   RECT 23.18 745.56 202.54 747.27 ;
   RECT 23.18 747.27 202.54 748.98 ;
   RECT 23.18 748.98 202.54 750.69 ;
   RECT 23.18 750.69 202.54 752.4 ;
   RECT 23.18 752.4 202.54 754.11 ;
   RECT 23.18 754.11 202.54 755.82 ;
   RECT 23.18 755.82 202.54 757.53 ;
   RECT 23.18 757.53 202.54 759.24 ;
   RECT 23.18 759.24 202.54 760.95 ;
   RECT 23.18 760.95 202.54 762.66 ;
   RECT 23.18 762.66 202.54 764.37 ;
   RECT 23.18 764.37 202.54 766.08 ;
   RECT 23.18 766.08 202.54 767.79 ;
   RECT 23.18 767.79 202.54 769.5 ;
   RECT 23.18 769.5 202.54 771.21 ;
   RECT 23.18 771.21 202.54 772.92 ;
   RECT 23.18 772.92 202.54 774.63 ;
   RECT 23.18 774.63 202.54 776.34 ;
   RECT 23.18 776.34 202.54 778.05 ;
   RECT 23.18 778.05 202.54 779.76 ;
   RECT 23.18 779.76 202.54 781.47 ;
   RECT 23.18 781.47 202.54 783.18 ;
   RECT 23.18 783.18 202.54 784.89 ;
   RECT 23.18 784.89 202.54 786.6 ;
   RECT 23.18 786.6 202.54 788.31 ;
   RECT 23.18 788.31 202.54 790.02 ;
   RECT 23.18 790.02 202.54 791.73 ;
   RECT 23.18 791.73 202.54 793.44 ;
   RECT 23.18 793.44 202.54 795.15 ;
   RECT 23.18 795.15 202.54 796.86 ;
   RECT 23.18 796.86 202.54 798.57 ;
   RECT 23.18 798.57 202.54 800.28 ;
   RECT 23.18 800.28 202.54 801.99 ;
   RECT 23.18 801.99 202.54 803.7 ;
   RECT 23.18 803.7 202.54 805.41 ;
   RECT 23.18 805.41 202.54 807.12 ;
   RECT 23.18 807.12 202.54 808.83 ;
   RECT 23.18 808.83 202.54 810.54 ;
   RECT 23.18 810.54 202.54 812.25 ;
   RECT 23.18 812.25 202.54 813.96 ;
   RECT 23.18 813.96 202.54 815.67 ;
   RECT 23.18 815.67 202.54 817.38 ;
   RECT 23.18 817.38 202.54 819.09 ;
   RECT 23.18 819.09 202.54 820.8 ;
   RECT 23.18 820.8 202.54 822.51 ;
   RECT 23.18 822.51 202.54 824.22 ;
   RECT 23.18 824.22 202.54 825.93 ;
   RECT 23.18 825.93 202.54 827.64 ;
   RECT 23.18 827.64 202.54 829.35 ;
   RECT 23.18 829.35 202.54 831.06 ;
   RECT 23.18 831.06 202.54 832.77 ;
   RECT 23.18 832.77 202.54 834.48 ;
   RECT 23.18 834.48 202.54 836.19 ;
   RECT 23.18 836.19 202.54 837.9 ;
   RECT 23.18 837.9 202.54 839.61 ;
   RECT 23.18 839.61 202.54 841.32 ;
  LAYER via2 ;
   RECT 23.18 0.0 202.54 1.71 ;
   RECT 23.18 1.71 202.54 3.42 ;
   RECT 23.18 3.42 202.54 5.13 ;
   RECT 23.18 5.13 202.54 6.84 ;
   RECT 23.18 6.84 202.54 8.55 ;
   RECT 23.18 8.55 202.54 10.26 ;
   RECT 23.18 10.26 202.54 11.97 ;
   RECT 23.18 11.97 202.54 13.68 ;
   RECT 23.18 13.68 202.54 15.39 ;
   RECT 23.18 15.39 202.54 17.1 ;
   RECT 23.18 17.1 202.54 18.81 ;
   RECT 23.18 18.81 202.54 20.52 ;
   RECT 23.18 20.52 202.54 22.23 ;
   RECT 23.18 22.23 202.54 23.94 ;
   RECT 23.18 23.94 202.54 25.65 ;
   RECT 23.18 25.65 202.54 27.36 ;
   RECT 23.18 27.36 202.54 29.07 ;
   RECT 23.18 29.07 202.54 30.78 ;
   RECT 23.18 30.78 202.54 32.49 ;
   RECT 23.18 32.49 202.54 34.2 ;
   RECT 23.18 34.2 202.54 35.91 ;
   RECT 23.18 35.91 202.54 37.62 ;
   RECT 23.18 37.62 202.54 39.33 ;
   RECT 23.18 39.33 202.54 41.04 ;
   RECT 23.18 41.04 202.54 42.75 ;
   RECT 23.18 42.75 202.54 44.46 ;
   RECT 23.18 44.46 202.54 46.17 ;
   RECT 23.18 46.17 202.54 47.88 ;
   RECT 23.18 47.88 202.54 49.59 ;
   RECT 23.18 49.59 202.54 51.3 ;
   RECT 23.18 51.3 202.54 53.01 ;
   RECT 23.18 53.01 202.54 54.72 ;
   RECT 23.18 54.72 202.54 56.43 ;
   RECT 23.18 56.43 202.54 58.14 ;
   RECT 23.18 58.14 202.54 59.85 ;
   RECT 23.18 59.85 202.54 61.56 ;
   RECT 23.18 61.56 202.54 63.27 ;
   RECT 23.18 63.27 202.54 64.98 ;
   RECT 23.18 64.98 202.54 66.69 ;
   RECT 23.18 66.69 202.54 68.4 ;
   RECT 23.18 68.4 202.54 70.11 ;
   RECT 23.18 70.11 202.54 71.82 ;
   RECT 23.18 71.82 202.54 73.53 ;
   RECT 23.18 73.53 202.54 75.24 ;
   RECT 23.18 75.24 202.54 76.95 ;
   RECT 23.18 76.95 202.54 78.66 ;
   RECT 23.18 78.66 202.54 80.37 ;
   RECT 23.18 80.37 202.54 82.08 ;
   RECT 23.18 82.08 202.54 83.79 ;
   RECT 23.18 83.79 202.54 85.5 ;
   RECT 23.18 85.5 202.54 87.21 ;
   RECT 23.18 87.21 202.54 88.92 ;
   RECT 23.18 88.92 202.54 90.63 ;
   RECT 23.18 90.63 202.54 92.34 ;
   RECT 23.18 92.34 202.54 94.05 ;
   RECT 23.18 94.05 202.54 95.76 ;
   RECT 23.18 95.76 202.54 97.47 ;
   RECT 23.18 97.47 202.54 99.18 ;
   RECT 23.18 99.18 202.54 100.89 ;
   RECT 23.18 100.89 202.54 102.6 ;
   RECT 23.18 102.6 202.54 104.31 ;
   RECT 23.18 104.31 202.54 106.02 ;
   RECT 23.18 106.02 202.54 107.73 ;
   RECT 23.18 107.73 202.54 109.44 ;
   RECT 23.18 109.44 202.54 111.15 ;
   RECT 23.18 111.15 202.54 112.86 ;
   RECT 23.18 112.86 202.54 114.57 ;
   RECT 23.18 114.57 202.54 116.28 ;
   RECT 23.18 116.28 202.54 117.99 ;
   RECT 23.18 117.99 202.54 119.7 ;
   RECT 23.18 119.7 202.54 121.41 ;
   RECT 23.18 121.41 202.54 123.12 ;
   RECT 23.18 123.12 202.54 124.83 ;
   RECT 23.18 124.83 202.54 126.54 ;
   RECT 23.18 126.54 202.54 128.25 ;
   RECT 23.18 128.25 202.54 129.96 ;
   RECT 23.18 129.96 202.54 131.67 ;
   RECT 23.18 131.67 202.54 133.38 ;
   RECT 23.18 133.38 202.54 135.09 ;
   RECT 23.18 135.09 202.54 136.8 ;
   RECT 23.18 136.8 202.54 138.51 ;
   RECT 23.18 138.51 202.54 140.22 ;
   RECT 23.18 140.22 202.54 141.93 ;
   RECT 23.18 141.93 202.54 143.64 ;
   RECT 23.18 143.64 202.54 145.35 ;
   RECT 23.18 145.35 202.54 147.06 ;
   RECT 23.18 147.06 202.54 148.77 ;
   RECT 23.18 148.77 202.54 150.48 ;
   RECT 23.18 150.48 202.54 152.19 ;
   RECT 23.18 152.19 202.54 153.9 ;
   RECT 23.18 153.9 202.54 155.61 ;
   RECT 23.18 155.61 202.54 157.32 ;
   RECT 23.18 157.32 202.54 159.03 ;
   RECT 23.18 159.03 202.54 160.74 ;
   RECT 23.18 160.74 202.54 162.45 ;
   RECT 23.18 162.45 202.54 164.16 ;
   RECT 23.18 164.16 202.54 165.87 ;
   RECT 23.18 165.87 202.54 167.58 ;
   RECT 23.18 167.58 202.54 169.29 ;
   RECT 23.18 169.29 202.54 171.0 ;
   RECT 23.18 171.0 202.54 172.71 ;
   RECT 23.18 172.71 202.54 174.42 ;
   RECT 23.18 174.42 202.54 176.13 ;
   RECT 23.18 176.13 202.54 177.84 ;
   RECT 23.18 177.84 202.54 179.55 ;
   RECT 23.18 179.55 202.54 181.26 ;
   RECT 23.18 181.26 202.54 182.97 ;
   RECT 23.18 182.97 202.54 184.68 ;
   RECT 23.18 184.68 202.54 186.39 ;
   RECT 23.18 186.39 202.54 188.1 ;
   RECT 23.18 188.1 202.54 189.81 ;
   RECT 23.18 189.81 202.54 191.52 ;
   RECT 23.18 191.52 202.54 193.23 ;
   RECT 23.18 193.23 202.54 194.94 ;
   RECT 23.18 194.94 202.54 196.65 ;
   RECT 23.18 196.65 202.54 198.36 ;
   RECT 23.18 198.36 202.54 200.07 ;
   RECT 23.18 200.07 202.54 201.78 ;
   RECT 23.18 201.78 202.54 203.49 ;
   RECT 23.18 203.49 202.54 205.2 ;
   RECT 23.18 205.2 202.54 206.91 ;
   RECT 23.18 206.91 202.54 208.62 ;
   RECT 23.18 208.62 202.54 210.33 ;
   RECT 23.18 210.33 202.54 212.04 ;
   RECT 23.18 212.04 202.54 213.75 ;
   RECT 23.18 213.75 202.54 215.46 ;
   RECT 23.18 215.46 202.54 217.17 ;
   RECT 23.18 217.17 202.54 218.88 ;
   RECT 23.18 218.88 202.54 220.59 ;
   RECT 23.18 220.59 202.54 222.3 ;
   RECT 23.18 222.3 202.54 224.01 ;
   RECT 23.18 224.01 202.54 225.72 ;
   RECT 23.18 225.72 202.54 227.43 ;
   RECT 23.18 227.43 202.54 229.14 ;
   RECT 23.18 229.14 202.54 230.85 ;
   RECT 23.18 230.85 202.54 232.56 ;
   RECT 23.18 232.56 202.54 234.27 ;
   RECT 23.18 234.27 202.54 235.98 ;
   RECT 23.18 235.98 202.54 237.69 ;
   RECT 23.18 237.69 202.54 239.4 ;
   RECT 23.18 239.4 202.54 241.11 ;
   RECT 23.18 241.11 202.54 242.82 ;
   RECT 23.18 242.82 202.54 244.53 ;
   RECT 23.18 244.53 202.54 246.24 ;
   RECT 23.18 246.24 202.54 247.95 ;
   RECT 23.18 247.95 202.54 249.66 ;
   RECT 23.18 249.66 202.54 251.37 ;
   RECT 23.18 251.37 202.54 253.08 ;
   RECT 23.18 253.08 202.54 254.79 ;
   RECT 23.18 254.79 202.54 256.5 ;
   RECT 23.18 256.5 202.54 258.21 ;
   RECT 23.18 258.21 202.54 259.92 ;
   RECT 23.18 259.92 202.54 261.63 ;
   RECT 23.18 261.63 202.54 263.34 ;
   RECT 23.18 263.34 202.54 265.05 ;
   RECT 23.18 265.05 202.54 266.76 ;
   RECT 23.18 266.76 202.54 268.47 ;
   RECT 23.18 268.47 202.54 270.18 ;
   RECT 23.18 270.18 202.54 271.89 ;
   RECT 23.18 271.89 202.54 273.6 ;
   RECT 23.18 273.6 202.54 275.31 ;
   RECT 23.18 275.31 202.54 277.02 ;
   RECT 23.18 277.02 202.54 278.73 ;
   RECT 23.18 278.73 202.54 280.44 ;
   RECT 23.18 280.44 202.54 282.15 ;
   RECT 23.18 282.15 202.54 283.86 ;
   RECT 23.18 283.86 202.54 285.57 ;
   RECT 23.18 285.57 202.54 287.28 ;
   RECT 23.18 287.28 202.54 288.99 ;
   RECT 23.18 288.99 202.54 290.7 ;
   RECT 23.18 290.7 202.54 292.41 ;
   RECT 23.18 292.41 202.54 294.12 ;
   RECT 23.18 294.12 202.54 295.83 ;
   RECT 23.18 295.83 202.54 297.54 ;
   RECT 23.18 297.54 202.54 299.25 ;
   RECT 23.18 299.25 202.54 300.96 ;
   RECT 23.18 300.96 202.54 302.67 ;
   RECT 23.18 302.67 202.54 304.38 ;
   RECT 23.18 304.38 202.54 306.09 ;
   RECT 23.18 306.09 202.54 307.8 ;
   RECT 23.18 307.8 202.54 309.51 ;
   RECT 23.18 309.51 202.54 311.22 ;
   RECT 23.18 311.22 202.54 312.93 ;
   RECT 23.18 312.93 202.54 314.64 ;
   RECT 23.18 314.64 202.54 316.35 ;
   RECT 23.18 316.35 202.54 318.06 ;
   RECT 23.18 318.06 202.54 319.77 ;
   RECT 23.18 319.77 202.54 321.48 ;
   RECT 23.18 321.48 202.54 323.19 ;
   RECT 23.18 323.19 202.54 324.9 ;
   RECT 23.18 324.9 202.54 326.61 ;
   RECT 23.18 326.61 202.54 328.32 ;
   RECT 23.18 328.32 202.54 330.03 ;
   RECT 23.18 330.03 202.54 331.74 ;
   RECT 23.18 331.74 202.54 333.45 ;
   RECT 23.18 333.45 202.54 335.16 ;
   RECT 23.18 335.16 202.54 336.87 ;
   RECT 23.18 336.87 202.54 338.58 ;
   RECT 23.18 338.58 202.54 340.29 ;
   RECT 23.18 340.29 202.54 342.0 ;
   RECT 23.18 342.0 202.54 343.71 ;
   RECT 23.18 343.71 202.54 345.42 ;
   RECT 23.18 345.42 202.54 347.13 ;
   RECT 23.18 347.13 202.54 348.84 ;
   RECT 23.18 348.84 202.54 350.55 ;
   RECT 23.18 350.55 202.54 352.26 ;
   RECT 23.18 352.26 202.54 353.97 ;
   RECT 23.18 353.97 202.54 355.68 ;
   RECT 23.18 355.68 202.54 357.39 ;
   RECT 23.18 357.39 202.54 359.1 ;
   RECT 23.18 359.1 202.54 360.81 ;
   RECT 23.18 360.81 202.54 362.52 ;
   RECT 23.18 362.52 202.54 364.23 ;
   RECT 23.18 364.23 202.54 365.94 ;
   RECT 23.18 365.94 202.54 367.65 ;
   RECT 23.18 367.65 202.54 369.36 ;
   RECT 23.18 369.36 202.54 371.07 ;
   RECT 23.18 371.07 202.54 372.78 ;
   RECT 23.18 372.78 202.54 374.49 ;
   RECT 23.18 374.49 202.54 376.2 ;
   RECT 23.18 376.2 202.54 377.91 ;
   RECT 23.18 377.91 202.54 379.62 ;
   RECT 23.18 379.62 202.54 381.33 ;
   RECT 23.18 381.33 202.54 383.04 ;
   RECT 23.18 383.04 202.54 384.75 ;
   RECT 23.18 384.75 202.54 386.46 ;
   RECT 23.18 386.46 202.54 388.17 ;
   RECT 23.18 388.17 202.54 389.88 ;
   RECT 23.18 389.88 202.54 391.59 ;
   RECT 23.18 391.59 202.54 393.3 ;
   RECT 23.18 393.3 202.54 395.01 ;
   RECT 23.18 395.01 202.54 396.72 ;
   RECT 23.18 396.72 202.54 398.43 ;
   RECT 23.18 398.43 202.54 400.14 ;
   RECT 23.18 400.14 202.54 401.85 ;
   RECT 0.0 401.85 202.54 403.56 ;
   RECT 0.0 403.56 202.54 405.27 ;
   RECT 0.0 405.27 202.54 406.98 ;
   RECT 0.0 406.98 202.54 408.69 ;
   RECT 0.0 408.69 202.54 410.4 ;
   RECT 0.0 410.4 202.54 412.11 ;
   RECT 0.0 412.11 202.54 413.82 ;
   RECT 0.0 413.82 202.54 415.53 ;
   RECT 0.0 415.53 202.54 417.24 ;
   RECT 0.0 417.24 202.54 418.95 ;
   RECT 0.0 418.95 202.54 420.66 ;
   RECT 0.0 420.66 202.54 422.37 ;
   RECT 0.0 422.37 202.54 424.08 ;
   RECT 0.0 424.08 202.54 425.79 ;
   RECT 0.0 425.79 202.54 427.5 ;
   RECT 0.0 427.5 202.54 429.21 ;
   RECT 0.0 429.21 202.54 430.92 ;
   RECT 23.18 430.92 202.54 432.63 ;
   RECT 23.18 432.63 202.54 434.34 ;
   RECT 23.18 434.34 202.54 436.05 ;
   RECT 23.18 436.05 202.54 437.76 ;
   RECT 23.18 437.76 202.54 439.47 ;
   RECT 23.18 439.47 202.54 441.18 ;
   RECT 23.18 441.18 202.54 442.89 ;
   RECT 23.18 442.89 202.54 444.6 ;
   RECT 23.18 444.6 202.54 446.31 ;
   RECT 23.18 446.31 202.54 448.02 ;
   RECT 23.18 448.02 202.54 449.73 ;
   RECT 23.18 449.73 202.54 451.44 ;
   RECT 23.18 451.44 202.54 453.15 ;
   RECT 23.18 453.15 202.54 454.86 ;
   RECT 23.18 454.86 202.54 456.57 ;
   RECT 23.18 456.57 202.54 458.28 ;
   RECT 23.18 458.28 202.54 459.99 ;
   RECT 23.18 459.99 202.54 461.7 ;
   RECT 23.18 461.7 202.54 463.41 ;
   RECT 23.18 463.41 202.54 465.12 ;
   RECT 23.18 465.12 202.54 466.83 ;
   RECT 23.18 466.83 202.54 468.54 ;
   RECT 23.18 468.54 202.54 470.25 ;
   RECT 23.18 470.25 202.54 471.96 ;
   RECT 23.18 471.96 202.54 473.67 ;
   RECT 23.18 473.67 202.54 475.38 ;
   RECT 23.18 475.38 202.54 477.09 ;
   RECT 23.18 477.09 202.54 478.8 ;
   RECT 23.18 478.8 202.54 480.51 ;
   RECT 23.18 480.51 202.54 482.22 ;
   RECT 23.18 482.22 202.54 483.93 ;
   RECT 23.18 483.93 202.54 485.64 ;
   RECT 23.18 485.64 202.54 487.35 ;
   RECT 23.18 487.35 202.54 489.06 ;
   RECT 23.18 489.06 202.54 490.77 ;
   RECT 23.18 490.77 202.54 492.48 ;
   RECT 23.18 492.48 202.54 494.19 ;
   RECT 23.18 494.19 202.54 495.9 ;
   RECT 23.18 495.9 202.54 497.61 ;
   RECT 23.18 497.61 202.54 499.32 ;
   RECT 23.18 499.32 202.54 501.03 ;
   RECT 23.18 501.03 202.54 502.74 ;
   RECT 23.18 502.74 202.54 504.45 ;
   RECT 23.18 504.45 202.54 506.16 ;
   RECT 23.18 506.16 202.54 507.87 ;
   RECT 23.18 507.87 202.54 509.58 ;
   RECT 23.18 509.58 202.54 511.29 ;
   RECT 23.18 511.29 202.54 513.0 ;
   RECT 23.18 513.0 202.54 514.71 ;
   RECT 23.18 514.71 202.54 516.42 ;
   RECT 23.18 516.42 202.54 518.13 ;
   RECT 23.18 518.13 202.54 519.84 ;
   RECT 23.18 519.84 202.54 521.55 ;
   RECT 23.18 521.55 202.54 523.26 ;
   RECT 23.18 523.26 202.54 524.97 ;
   RECT 23.18 524.97 202.54 526.68 ;
   RECT 23.18 526.68 202.54 528.39 ;
   RECT 23.18 528.39 202.54 530.1 ;
   RECT 23.18 530.1 202.54 531.81 ;
   RECT 23.18 531.81 202.54 533.52 ;
   RECT 23.18 533.52 202.54 535.23 ;
   RECT 23.18 535.23 202.54 536.94 ;
   RECT 23.18 536.94 202.54 538.65 ;
   RECT 23.18 538.65 202.54 540.36 ;
   RECT 23.18 540.36 202.54 542.07 ;
   RECT 23.18 542.07 202.54 543.78 ;
   RECT 23.18 543.78 202.54 545.49 ;
   RECT 23.18 545.49 202.54 547.2 ;
   RECT 23.18 547.2 202.54 548.91 ;
   RECT 23.18 548.91 202.54 550.62 ;
   RECT 23.18 550.62 202.54 552.33 ;
   RECT 23.18 552.33 202.54 554.04 ;
   RECT 23.18 554.04 202.54 555.75 ;
   RECT 23.18 555.75 202.54 557.46 ;
   RECT 23.18 557.46 202.54 559.17 ;
   RECT 23.18 559.17 202.54 560.88 ;
   RECT 23.18 560.88 202.54 562.59 ;
   RECT 23.18 562.59 202.54 564.3 ;
   RECT 23.18 564.3 202.54 566.01 ;
   RECT 23.18 566.01 202.54 567.72 ;
   RECT 23.18 567.72 202.54 569.43 ;
   RECT 23.18 569.43 202.54 571.14 ;
   RECT 23.18 571.14 202.54 572.85 ;
   RECT 23.18 572.85 202.54 574.56 ;
   RECT 23.18 574.56 202.54 576.27 ;
   RECT 23.18 576.27 202.54 577.98 ;
   RECT 23.18 577.98 202.54 579.69 ;
   RECT 23.18 579.69 202.54 581.4 ;
   RECT 23.18 581.4 202.54 583.11 ;
   RECT 23.18 583.11 202.54 584.82 ;
   RECT 23.18 584.82 202.54 586.53 ;
   RECT 23.18 586.53 202.54 588.24 ;
   RECT 23.18 588.24 202.54 589.95 ;
   RECT 23.18 589.95 202.54 591.66 ;
   RECT 23.18 591.66 202.54 593.37 ;
   RECT 23.18 593.37 202.54 595.08 ;
   RECT 23.18 595.08 202.54 596.79 ;
   RECT 23.18 596.79 202.54 598.5 ;
   RECT 23.18 598.5 202.54 600.21 ;
   RECT 23.18 600.21 202.54 601.92 ;
   RECT 23.18 601.92 202.54 603.63 ;
   RECT 23.18 603.63 202.54 605.34 ;
   RECT 23.18 605.34 202.54 607.05 ;
   RECT 23.18 607.05 202.54 608.76 ;
   RECT 23.18 608.76 202.54 610.47 ;
   RECT 23.18 610.47 202.54 612.18 ;
   RECT 23.18 612.18 202.54 613.89 ;
   RECT 23.18 613.89 202.54 615.6 ;
   RECT 23.18 615.6 202.54 617.31 ;
   RECT 23.18 617.31 202.54 619.02 ;
   RECT 23.18 619.02 202.54 620.73 ;
   RECT 23.18 620.73 202.54 622.44 ;
   RECT 23.18 622.44 202.54 624.15 ;
   RECT 23.18 624.15 202.54 625.86 ;
   RECT 23.18 625.86 202.54 627.57 ;
   RECT 23.18 627.57 202.54 629.28 ;
   RECT 23.18 629.28 202.54 630.99 ;
   RECT 23.18 630.99 202.54 632.7 ;
   RECT 23.18 632.7 202.54 634.41 ;
   RECT 23.18 634.41 202.54 636.12 ;
   RECT 23.18 636.12 202.54 637.83 ;
   RECT 23.18 637.83 202.54 639.54 ;
   RECT 23.18 639.54 202.54 641.25 ;
   RECT 23.18 641.25 202.54 642.96 ;
   RECT 23.18 642.96 202.54 644.67 ;
   RECT 23.18 644.67 202.54 646.38 ;
   RECT 23.18 646.38 202.54 648.09 ;
   RECT 23.18 648.09 202.54 649.8 ;
   RECT 23.18 649.8 202.54 651.51 ;
   RECT 23.18 651.51 202.54 653.22 ;
   RECT 23.18 653.22 202.54 654.93 ;
   RECT 23.18 654.93 202.54 656.64 ;
   RECT 23.18 656.64 202.54 658.35 ;
   RECT 23.18 658.35 202.54 660.06 ;
   RECT 23.18 660.06 202.54 661.77 ;
   RECT 23.18 661.77 202.54 663.48 ;
   RECT 23.18 663.48 202.54 665.19 ;
   RECT 23.18 665.19 202.54 666.9 ;
   RECT 23.18 666.9 202.54 668.61 ;
   RECT 23.18 668.61 202.54 670.32 ;
   RECT 23.18 670.32 202.54 672.03 ;
   RECT 23.18 672.03 202.54 673.74 ;
   RECT 23.18 673.74 202.54 675.45 ;
   RECT 23.18 675.45 202.54 677.16 ;
   RECT 23.18 677.16 202.54 678.87 ;
   RECT 23.18 678.87 202.54 680.58 ;
   RECT 23.18 680.58 202.54 682.29 ;
   RECT 23.18 682.29 202.54 684.0 ;
   RECT 23.18 684.0 202.54 685.71 ;
   RECT 23.18 685.71 202.54 687.42 ;
   RECT 23.18 687.42 202.54 689.13 ;
   RECT 23.18 689.13 202.54 690.84 ;
   RECT 23.18 690.84 202.54 692.55 ;
   RECT 23.18 692.55 202.54 694.26 ;
   RECT 23.18 694.26 202.54 695.97 ;
   RECT 23.18 695.97 202.54 697.68 ;
   RECT 23.18 697.68 202.54 699.39 ;
   RECT 23.18 699.39 202.54 701.1 ;
   RECT 23.18 701.1 202.54 702.81 ;
   RECT 23.18 702.81 202.54 704.52 ;
   RECT 23.18 704.52 202.54 706.23 ;
   RECT 23.18 706.23 202.54 707.94 ;
   RECT 23.18 707.94 202.54 709.65 ;
   RECT 23.18 709.65 202.54 711.36 ;
   RECT 23.18 711.36 202.54 713.07 ;
   RECT 23.18 713.07 202.54 714.78 ;
   RECT 23.18 714.78 202.54 716.49 ;
   RECT 23.18 716.49 202.54 718.2 ;
   RECT 23.18 718.2 202.54 719.91 ;
   RECT 23.18 719.91 202.54 721.62 ;
   RECT 23.18 721.62 202.54 723.33 ;
   RECT 23.18 723.33 202.54 725.04 ;
   RECT 23.18 725.04 202.54 726.75 ;
   RECT 23.18 726.75 202.54 728.46 ;
   RECT 23.18 728.46 202.54 730.17 ;
   RECT 23.18 730.17 202.54 731.88 ;
   RECT 23.18 731.88 202.54 733.59 ;
   RECT 23.18 733.59 202.54 735.3 ;
   RECT 23.18 735.3 202.54 737.01 ;
   RECT 23.18 737.01 202.54 738.72 ;
   RECT 23.18 738.72 202.54 740.43 ;
   RECT 23.18 740.43 202.54 742.14 ;
   RECT 23.18 742.14 202.54 743.85 ;
   RECT 23.18 743.85 202.54 745.56 ;
   RECT 23.18 745.56 202.54 747.27 ;
   RECT 23.18 747.27 202.54 748.98 ;
   RECT 23.18 748.98 202.54 750.69 ;
   RECT 23.18 750.69 202.54 752.4 ;
   RECT 23.18 752.4 202.54 754.11 ;
   RECT 23.18 754.11 202.54 755.82 ;
   RECT 23.18 755.82 202.54 757.53 ;
   RECT 23.18 757.53 202.54 759.24 ;
   RECT 23.18 759.24 202.54 760.95 ;
   RECT 23.18 760.95 202.54 762.66 ;
   RECT 23.18 762.66 202.54 764.37 ;
   RECT 23.18 764.37 202.54 766.08 ;
   RECT 23.18 766.08 202.54 767.79 ;
   RECT 23.18 767.79 202.54 769.5 ;
   RECT 23.18 769.5 202.54 771.21 ;
   RECT 23.18 771.21 202.54 772.92 ;
   RECT 23.18 772.92 202.54 774.63 ;
   RECT 23.18 774.63 202.54 776.34 ;
   RECT 23.18 776.34 202.54 778.05 ;
   RECT 23.18 778.05 202.54 779.76 ;
   RECT 23.18 779.76 202.54 781.47 ;
   RECT 23.18 781.47 202.54 783.18 ;
   RECT 23.18 783.18 202.54 784.89 ;
   RECT 23.18 784.89 202.54 786.6 ;
   RECT 23.18 786.6 202.54 788.31 ;
   RECT 23.18 788.31 202.54 790.02 ;
   RECT 23.18 790.02 202.54 791.73 ;
   RECT 23.18 791.73 202.54 793.44 ;
   RECT 23.18 793.44 202.54 795.15 ;
   RECT 23.18 795.15 202.54 796.86 ;
   RECT 23.18 796.86 202.54 798.57 ;
   RECT 23.18 798.57 202.54 800.28 ;
   RECT 23.18 800.28 202.54 801.99 ;
   RECT 23.18 801.99 202.54 803.7 ;
   RECT 23.18 803.7 202.54 805.41 ;
   RECT 23.18 805.41 202.54 807.12 ;
   RECT 23.18 807.12 202.54 808.83 ;
   RECT 23.18 808.83 202.54 810.54 ;
   RECT 23.18 810.54 202.54 812.25 ;
   RECT 23.18 812.25 202.54 813.96 ;
   RECT 23.18 813.96 202.54 815.67 ;
   RECT 23.18 815.67 202.54 817.38 ;
   RECT 23.18 817.38 202.54 819.09 ;
   RECT 23.18 819.09 202.54 820.8 ;
   RECT 23.18 820.8 202.54 822.51 ;
   RECT 23.18 822.51 202.54 824.22 ;
   RECT 23.18 824.22 202.54 825.93 ;
   RECT 23.18 825.93 202.54 827.64 ;
   RECT 23.18 827.64 202.54 829.35 ;
   RECT 23.18 829.35 202.54 831.06 ;
   RECT 23.18 831.06 202.54 832.77 ;
   RECT 23.18 832.77 202.54 834.48 ;
   RECT 23.18 834.48 202.54 836.19 ;
   RECT 23.18 836.19 202.54 837.9 ;
   RECT 23.18 837.9 202.54 839.61 ;
   RECT 23.18 839.61 202.54 841.32 ;
  LAYER metal3 ;
   RECT 23.18 0.0 202.54 1.71 ;
   RECT 23.18 1.71 202.54 3.42 ;
   RECT 23.18 3.42 202.54 5.13 ;
   RECT 23.18 5.13 202.54 6.84 ;
   RECT 23.18 6.84 202.54 8.55 ;
   RECT 23.18 8.55 202.54 10.26 ;
   RECT 23.18 10.26 202.54 11.97 ;
   RECT 23.18 11.97 202.54 13.68 ;
   RECT 23.18 13.68 202.54 15.39 ;
   RECT 23.18 15.39 202.54 17.1 ;
   RECT 23.18 17.1 202.54 18.81 ;
   RECT 23.18 18.81 202.54 20.52 ;
   RECT 23.18 20.52 202.54 22.23 ;
   RECT 23.18 22.23 202.54 23.94 ;
   RECT 23.18 23.94 202.54 25.65 ;
   RECT 23.18 25.65 202.54 27.36 ;
   RECT 23.18 27.36 202.54 29.07 ;
   RECT 23.18 29.07 202.54 30.78 ;
   RECT 23.18 30.78 202.54 32.49 ;
   RECT 23.18 32.49 202.54 34.2 ;
   RECT 23.18 34.2 202.54 35.91 ;
   RECT 23.18 35.91 202.54 37.62 ;
   RECT 23.18 37.62 202.54 39.33 ;
   RECT 23.18 39.33 202.54 41.04 ;
   RECT 23.18 41.04 202.54 42.75 ;
   RECT 23.18 42.75 202.54 44.46 ;
   RECT 23.18 44.46 202.54 46.17 ;
   RECT 23.18 46.17 202.54 47.88 ;
   RECT 23.18 47.88 202.54 49.59 ;
   RECT 23.18 49.59 202.54 51.3 ;
   RECT 23.18 51.3 202.54 53.01 ;
   RECT 23.18 53.01 202.54 54.72 ;
   RECT 23.18 54.72 202.54 56.43 ;
   RECT 23.18 56.43 202.54 58.14 ;
   RECT 23.18 58.14 202.54 59.85 ;
   RECT 23.18 59.85 202.54 61.56 ;
   RECT 23.18 61.56 202.54 63.27 ;
   RECT 23.18 63.27 202.54 64.98 ;
   RECT 23.18 64.98 202.54 66.69 ;
   RECT 23.18 66.69 202.54 68.4 ;
   RECT 23.18 68.4 202.54 70.11 ;
   RECT 23.18 70.11 202.54 71.82 ;
   RECT 23.18 71.82 202.54 73.53 ;
   RECT 23.18 73.53 202.54 75.24 ;
   RECT 23.18 75.24 202.54 76.95 ;
   RECT 23.18 76.95 202.54 78.66 ;
   RECT 23.18 78.66 202.54 80.37 ;
   RECT 23.18 80.37 202.54 82.08 ;
   RECT 23.18 82.08 202.54 83.79 ;
   RECT 23.18 83.79 202.54 85.5 ;
   RECT 23.18 85.5 202.54 87.21 ;
   RECT 23.18 87.21 202.54 88.92 ;
   RECT 23.18 88.92 202.54 90.63 ;
   RECT 23.18 90.63 202.54 92.34 ;
   RECT 23.18 92.34 202.54 94.05 ;
   RECT 23.18 94.05 202.54 95.76 ;
   RECT 23.18 95.76 202.54 97.47 ;
   RECT 23.18 97.47 202.54 99.18 ;
   RECT 23.18 99.18 202.54 100.89 ;
   RECT 23.18 100.89 202.54 102.6 ;
   RECT 23.18 102.6 202.54 104.31 ;
   RECT 23.18 104.31 202.54 106.02 ;
   RECT 23.18 106.02 202.54 107.73 ;
   RECT 23.18 107.73 202.54 109.44 ;
   RECT 23.18 109.44 202.54 111.15 ;
   RECT 23.18 111.15 202.54 112.86 ;
   RECT 23.18 112.86 202.54 114.57 ;
   RECT 23.18 114.57 202.54 116.28 ;
   RECT 23.18 116.28 202.54 117.99 ;
   RECT 23.18 117.99 202.54 119.7 ;
   RECT 23.18 119.7 202.54 121.41 ;
   RECT 23.18 121.41 202.54 123.12 ;
   RECT 23.18 123.12 202.54 124.83 ;
   RECT 23.18 124.83 202.54 126.54 ;
   RECT 23.18 126.54 202.54 128.25 ;
   RECT 23.18 128.25 202.54 129.96 ;
   RECT 23.18 129.96 202.54 131.67 ;
   RECT 23.18 131.67 202.54 133.38 ;
   RECT 23.18 133.38 202.54 135.09 ;
   RECT 23.18 135.09 202.54 136.8 ;
   RECT 23.18 136.8 202.54 138.51 ;
   RECT 23.18 138.51 202.54 140.22 ;
   RECT 23.18 140.22 202.54 141.93 ;
   RECT 23.18 141.93 202.54 143.64 ;
   RECT 23.18 143.64 202.54 145.35 ;
   RECT 23.18 145.35 202.54 147.06 ;
   RECT 23.18 147.06 202.54 148.77 ;
   RECT 23.18 148.77 202.54 150.48 ;
   RECT 23.18 150.48 202.54 152.19 ;
   RECT 23.18 152.19 202.54 153.9 ;
   RECT 23.18 153.9 202.54 155.61 ;
   RECT 23.18 155.61 202.54 157.32 ;
   RECT 23.18 157.32 202.54 159.03 ;
   RECT 23.18 159.03 202.54 160.74 ;
   RECT 23.18 160.74 202.54 162.45 ;
   RECT 23.18 162.45 202.54 164.16 ;
   RECT 23.18 164.16 202.54 165.87 ;
   RECT 23.18 165.87 202.54 167.58 ;
   RECT 23.18 167.58 202.54 169.29 ;
   RECT 23.18 169.29 202.54 171.0 ;
   RECT 23.18 171.0 202.54 172.71 ;
   RECT 23.18 172.71 202.54 174.42 ;
   RECT 23.18 174.42 202.54 176.13 ;
   RECT 23.18 176.13 202.54 177.84 ;
   RECT 23.18 177.84 202.54 179.55 ;
   RECT 23.18 179.55 202.54 181.26 ;
   RECT 23.18 181.26 202.54 182.97 ;
   RECT 23.18 182.97 202.54 184.68 ;
   RECT 23.18 184.68 202.54 186.39 ;
   RECT 23.18 186.39 202.54 188.1 ;
   RECT 23.18 188.1 202.54 189.81 ;
   RECT 23.18 189.81 202.54 191.52 ;
   RECT 23.18 191.52 202.54 193.23 ;
   RECT 23.18 193.23 202.54 194.94 ;
   RECT 23.18 194.94 202.54 196.65 ;
   RECT 23.18 196.65 202.54 198.36 ;
   RECT 23.18 198.36 202.54 200.07 ;
   RECT 23.18 200.07 202.54 201.78 ;
   RECT 23.18 201.78 202.54 203.49 ;
   RECT 23.18 203.49 202.54 205.2 ;
   RECT 23.18 205.2 202.54 206.91 ;
   RECT 23.18 206.91 202.54 208.62 ;
   RECT 23.18 208.62 202.54 210.33 ;
   RECT 23.18 210.33 202.54 212.04 ;
   RECT 23.18 212.04 202.54 213.75 ;
   RECT 23.18 213.75 202.54 215.46 ;
   RECT 23.18 215.46 202.54 217.17 ;
   RECT 23.18 217.17 202.54 218.88 ;
   RECT 23.18 218.88 202.54 220.59 ;
   RECT 23.18 220.59 202.54 222.3 ;
   RECT 23.18 222.3 202.54 224.01 ;
   RECT 23.18 224.01 202.54 225.72 ;
   RECT 23.18 225.72 202.54 227.43 ;
   RECT 23.18 227.43 202.54 229.14 ;
   RECT 23.18 229.14 202.54 230.85 ;
   RECT 23.18 230.85 202.54 232.56 ;
   RECT 23.18 232.56 202.54 234.27 ;
   RECT 23.18 234.27 202.54 235.98 ;
   RECT 23.18 235.98 202.54 237.69 ;
   RECT 23.18 237.69 202.54 239.4 ;
   RECT 23.18 239.4 202.54 241.11 ;
   RECT 23.18 241.11 202.54 242.82 ;
   RECT 23.18 242.82 202.54 244.53 ;
   RECT 23.18 244.53 202.54 246.24 ;
   RECT 23.18 246.24 202.54 247.95 ;
   RECT 23.18 247.95 202.54 249.66 ;
   RECT 23.18 249.66 202.54 251.37 ;
   RECT 23.18 251.37 202.54 253.08 ;
   RECT 23.18 253.08 202.54 254.79 ;
   RECT 23.18 254.79 202.54 256.5 ;
   RECT 23.18 256.5 202.54 258.21 ;
   RECT 23.18 258.21 202.54 259.92 ;
   RECT 23.18 259.92 202.54 261.63 ;
   RECT 23.18 261.63 202.54 263.34 ;
   RECT 23.18 263.34 202.54 265.05 ;
   RECT 23.18 265.05 202.54 266.76 ;
   RECT 23.18 266.76 202.54 268.47 ;
   RECT 23.18 268.47 202.54 270.18 ;
   RECT 23.18 270.18 202.54 271.89 ;
   RECT 23.18 271.89 202.54 273.6 ;
   RECT 23.18 273.6 202.54 275.31 ;
   RECT 23.18 275.31 202.54 277.02 ;
   RECT 23.18 277.02 202.54 278.73 ;
   RECT 23.18 278.73 202.54 280.44 ;
   RECT 23.18 280.44 202.54 282.15 ;
   RECT 23.18 282.15 202.54 283.86 ;
   RECT 23.18 283.86 202.54 285.57 ;
   RECT 23.18 285.57 202.54 287.28 ;
   RECT 23.18 287.28 202.54 288.99 ;
   RECT 23.18 288.99 202.54 290.7 ;
   RECT 23.18 290.7 202.54 292.41 ;
   RECT 23.18 292.41 202.54 294.12 ;
   RECT 23.18 294.12 202.54 295.83 ;
   RECT 23.18 295.83 202.54 297.54 ;
   RECT 23.18 297.54 202.54 299.25 ;
   RECT 23.18 299.25 202.54 300.96 ;
   RECT 23.18 300.96 202.54 302.67 ;
   RECT 23.18 302.67 202.54 304.38 ;
   RECT 23.18 304.38 202.54 306.09 ;
   RECT 23.18 306.09 202.54 307.8 ;
   RECT 23.18 307.8 202.54 309.51 ;
   RECT 23.18 309.51 202.54 311.22 ;
   RECT 23.18 311.22 202.54 312.93 ;
   RECT 23.18 312.93 202.54 314.64 ;
   RECT 23.18 314.64 202.54 316.35 ;
   RECT 23.18 316.35 202.54 318.06 ;
   RECT 23.18 318.06 202.54 319.77 ;
   RECT 23.18 319.77 202.54 321.48 ;
   RECT 23.18 321.48 202.54 323.19 ;
   RECT 23.18 323.19 202.54 324.9 ;
   RECT 23.18 324.9 202.54 326.61 ;
   RECT 23.18 326.61 202.54 328.32 ;
   RECT 23.18 328.32 202.54 330.03 ;
   RECT 23.18 330.03 202.54 331.74 ;
   RECT 23.18 331.74 202.54 333.45 ;
   RECT 23.18 333.45 202.54 335.16 ;
   RECT 23.18 335.16 202.54 336.87 ;
   RECT 23.18 336.87 202.54 338.58 ;
   RECT 23.18 338.58 202.54 340.29 ;
   RECT 23.18 340.29 202.54 342.0 ;
   RECT 23.18 342.0 202.54 343.71 ;
   RECT 23.18 343.71 202.54 345.42 ;
   RECT 23.18 345.42 202.54 347.13 ;
   RECT 23.18 347.13 202.54 348.84 ;
   RECT 23.18 348.84 202.54 350.55 ;
   RECT 23.18 350.55 202.54 352.26 ;
   RECT 23.18 352.26 202.54 353.97 ;
   RECT 23.18 353.97 202.54 355.68 ;
   RECT 23.18 355.68 202.54 357.39 ;
   RECT 23.18 357.39 202.54 359.1 ;
   RECT 23.18 359.1 202.54 360.81 ;
   RECT 23.18 360.81 202.54 362.52 ;
   RECT 23.18 362.52 202.54 364.23 ;
   RECT 23.18 364.23 202.54 365.94 ;
   RECT 23.18 365.94 202.54 367.65 ;
   RECT 23.18 367.65 202.54 369.36 ;
   RECT 23.18 369.36 202.54 371.07 ;
   RECT 23.18 371.07 202.54 372.78 ;
   RECT 23.18 372.78 202.54 374.49 ;
   RECT 23.18 374.49 202.54 376.2 ;
   RECT 23.18 376.2 202.54 377.91 ;
   RECT 23.18 377.91 202.54 379.62 ;
   RECT 23.18 379.62 202.54 381.33 ;
   RECT 23.18 381.33 202.54 383.04 ;
   RECT 23.18 383.04 202.54 384.75 ;
   RECT 23.18 384.75 202.54 386.46 ;
   RECT 23.18 386.46 202.54 388.17 ;
   RECT 23.18 388.17 202.54 389.88 ;
   RECT 23.18 389.88 202.54 391.59 ;
   RECT 23.18 391.59 202.54 393.3 ;
   RECT 23.18 393.3 202.54 395.01 ;
   RECT 23.18 395.01 202.54 396.72 ;
   RECT 23.18 396.72 202.54 398.43 ;
   RECT 23.18 398.43 202.54 400.14 ;
   RECT 23.18 400.14 202.54 401.85 ;
   RECT 0.0 401.85 202.54 403.56 ;
   RECT 0.0 403.56 202.54 405.27 ;
   RECT 0.0 405.27 202.54 406.98 ;
   RECT 0.0 406.98 202.54 408.69 ;
   RECT 0.0 408.69 202.54 410.4 ;
   RECT 0.0 410.4 202.54 412.11 ;
   RECT 0.0 412.11 202.54 413.82 ;
   RECT 0.0 413.82 202.54 415.53 ;
   RECT 0.0 415.53 202.54 417.24 ;
   RECT 0.0 417.24 202.54 418.95 ;
   RECT 0.0 418.95 202.54 420.66 ;
   RECT 0.0 420.66 202.54 422.37 ;
   RECT 0.0 422.37 202.54 424.08 ;
   RECT 0.0 424.08 202.54 425.79 ;
   RECT 0.0 425.79 202.54 427.5 ;
   RECT 0.0 427.5 202.54 429.21 ;
   RECT 0.0 429.21 202.54 430.92 ;
   RECT 23.18 430.92 202.54 432.63 ;
   RECT 23.18 432.63 202.54 434.34 ;
   RECT 23.18 434.34 202.54 436.05 ;
   RECT 23.18 436.05 202.54 437.76 ;
   RECT 23.18 437.76 202.54 439.47 ;
   RECT 23.18 439.47 202.54 441.18 ;
   RECT 23.18 441.18 202.54 442.89 ;
   RECT 23.18 442.89 202.54 444.6 ;
   RECT 23.18 444.6 202.54 446.31 ;
   RECT 23.18 446.31 202.54 448.02 ;
   RECT 23.18 448.02 202.54 449.73 ;
   RECT 23.18 449.73 202.54 451.44 ;
   RECT 23.18 451.44 202.54 453.15 ;
   RECT 23.18 453.15 202.54 454.86 ;
   RECT 23.18 454.86 202.54 456.57 ;
   RECT 23.18 456.57 202.54 458.28 ;
   RECT 23.18 458.28 202.54 459.99 ;
   RECT 23.18 459.99 202.54 461.7 ;
   RECT 23.18 461.7 202.54 463.41 ;
   RECT 23.18 463.41 202.54 465.12 ;
   RECT 23.18 465.12 202.54 466.83 ;
   RECT 23.18 466.83 202.54 468.54 ;
   RECT 23.18 468.54 202.54 470.25 ;
   RECT 23.18 470.25 202.54 471.96 ;
   RECT 23.18 471.96 202.54 473.67 ;
   RECT 23.18 473.67 202.54 475.38 ;
   RECT 23.18 475.38 202.54 477.09 ;
   RECT 23.18 477.09 202.54 478.8 ;
   RECT 23.18 478.8 202.54 480.51 ;
   RECT 23.18 480.51 202.54 482.22 ;
   RECT 23.18 482.22 202.54 483.93 ;
   RECT 23.18 483.93 202.54 485.64 ;
   RECT 23.18 485.64 202.54 487.35 ;
   RECT 23.18 487.35 202.54 489.06 ;
   RECT 23.18 489.06 202.54 490.77 ;
   RECT 23.18 490.77 202.54 492.48 ;
   RECT 23.18 492.48 202.54 494.19 ;
   RECT 23.18 494.19 202.54 495.9 ;
   RECT 23.18 495.9 202.54 497.61 ;
   RECT 23.18 497.61 202.54 499.32 ;
   RECT 23.18 499.32 202.54 501.03 ;
   RECT 23.18 501.03 202.54 502.74 ;
   RECT 23.18 502.74 202.54 504.45 ;
   RECT 23.18 504.45 202.54 506.16 ;
   RECT 23.18 506.16 202.54 507.87 ;
   RECT 23.18 507.87 202.54 509.58 ;
   RECT 23.18 509.58 202.54 511.29 ;
   RECT 23.18 511.29 202.54 513.0 ;
   RECT 23.18 513.0 202.54 514.71 ;
   RECT 23.18 514.71 202.54 516.42 ;
   RECT 23.18 516.42 202.54 518.13 ;
   RECT 23.18 518.13 202.54 519.84 ;
   RECT 23.18 519.84 202.54 521.55 ;
   RECT 23.18 521.55 202.54 523.26 ;
   RECT 23.18 523.26 202.54 524.97 ;
   RECT 23.18 524.97 202.54 526.68 ;
   RECT 23.18 526.68 202.54 528.39 ;
   RECT 23.18 528.39 202.54 530.1 ;
   RECT 23.18 530.1 202.54 531.81 ;
   RECT 23.18 531.81 202.54 533.52 ;
   RECT 23.18 533.52 202.54 535.23 ;
   RECT 23.18 535.23 202.54 536.94 ;
   RECT 23.18 536.94 202.54 538.65 ;
   RECT 23.18 538.65 202.54 540.36 ;
   RECT 23.18 540.36 202.54 542.07 ;
   RECT 23.18 542.07 202.54 543.78 ;
   RECT 23.18 543.78 202.54 545.49 ;
   RECT 23.18 545.49 202.54 547.2 ;
   RECT 23.18 547.2 202.54 548.91 ;
   RECT 23.18 548.91 202.54 550.62 ;
   RECT 23.18 550.62 202.54 552.33 ;
   RECT 23.18 552.33 202.54 554.04 ;
   RECT 23.18 554.04 202.54 555.75 ;
   RECT 23.18 555.75 202.54 557.46 ;
   RECT 23.18 557.46 202.54 559.17 ;
   RECT 23.18 559.17 202.54 560.88 ;
   RECT 23.18 560.88 202.54 562.59 ;
   RECT 23.18 562.59 202.54 564.3 ;
   RECT 23.18 564.3 202.54 566.01 ;
   RECT 23.18 566.01 202.54 567.72 ;
   RECT 23.18 567.72 202.54 569.43 ;
   RECT 23.18 569.43 202.54 571.14 ;
   RECT 23.18 571.14 202.54 572.85 ;
   RECT 23.18 572.85 202.54 574.56 ;
   RECT 23.18 574.56 202.54 576.27 ;
   RECT 23.18 576.27 202.54 577.98 ;
   RECT 23.18 577.98 202.54 579.69 ;
   RECT 23.18 579.69 202.54 581.4 ;
   RECT 23.18 581.4 202.54 583.11 ;
   RECT 23.18 583.11 202.54 584.82 ;
   RECT 23.18 584.82 202.54 586.53 ;
   RECT 23.18 586.53 202.54 588.24 ;
   RECT 23.18 588.24 202.54 589.95 ;
   RECT 23.18 589.95 202.54 591.66 ;
   RECT 23.18 591.66 202.54 593.37 ;
   RECT 23.18 593.37 202.54 595.08 ;
   RECT 23.18 595.08 202.54 596.79 ;
   RECT 23.18 596.79 202.54 598.5 ;
   RECT 23.18 598.5 202.54 600.21 ;
   RECT 23.18 600.21 202.54 601.92 ;
   RECT 23.18 601.92 202.54 603.63 ;
   RECT 23.18 603.63 202.54 605.34 ;
   RECT 23.18 605.34 202.54 607.05 ;
   RECT 23.18 607.05 202.54 608.76 ;
   RECT 23.18 608.76 202.54 610.47 ;
   RECT 23.18 610.47 202.54 612.18 ;
   RECT 23.18 612.18 202.54 613.89 ;
   RECT 23.18 613.89 202.54 615.6 ;
   RECT 23.18 615.6 202.54 617.31 ;
   RECT 23.18 617.31 202.54 619.02 ;
   RECT 23.18 619.02 202.54 620.73 ;
   RECT 23.18 620.73 202.54 622.44 ;
   RECT 23.18 622.44 202.54 624.15 ;
   RECT 23.18 624.15 202.54 625.86 ;
   RECT 23.18 625.86 202.54 627.57 ;
   RECT 23.18 627.57 202.54 629.28 ;
   RECT 23.18 629.28 202.54 630.99 ;
   RECT 23.18 630.99 202.54 632.7 ;
   RECT 23.18 632.7 202.54 634.41 ;
   RECT 23.18 634.41 202.54 636.12 ;
   RECT 23.18 636.12 202.54 637.83 ;
   RECT 23.18 637.83 202.54 639.54 ;
   RECT 23.18 639.54 202.54 641.25 ;
   RECT 23.18 641.25 202.54 642.96 ;
   RECT 23.18 642.96 202.54 644.67 ;
   RECT 23.18 644.67 202.54 646.38 ;
   RECT 23.18 646.38 202.54 648.09 ;
   RECT 23.18 648.09 202.54 649.8 ;
   RECT 23.18 649.8 202.54 651.51 ;
   RECT 23.18 651.51 202.54 653.22 ;
   RECT 23.18 653.22 202.54 654.93 ;
   RECT 23.18 654.93 202.54 656.64 ;
   RECT 23.18 656.64 202.54 658.35 ;
   RECT 23.18 658.35 202.54 660.06 ;
   RECT 23.18 660.06 202.54 661.77 ;
   RECT 23.18 661.77 202.54 663.48 ;
   RECT 23.18 663.48 202.54 665.19 ;
   RECT 23.18 665.19 202.54 666.9 ;
   RECT 23.18 666.9 202.54 668.61 ;
   RECT 23.18 668.61 202.54 670.32 ;
   RECT 23.18 670.32 202.54 672.03 ;
   RECT 23.18 672.03 202.54 673.74 ;
   RECT 23.18 673.74 202.54 675.45 ;
   RECT 23.18 675.45 202.54 677.16 ;
   RECT 23.18 677.16 202.54 678.87 ;
   RECT 23.18 678.87 202.54 680.58 ;
   RECT 23.18 680.58 202.54 682.29 ;
   RECT 23.18 682.29 202.54 684.0 ;
   RECT 23.18 684.0 202.54 685.71 ;
   RECT 23.18 685.71 202.54 687.42 ;
   RECT 23.18 687.42 202.54 689.13 ;
   RECT 23.18 689.13 202.54 690.84 ;
   RECT 23.18 690.84 202.54 692.55 ;
   RECT 23.18 692.55 202.54 694.26 ;
   RECT 23.18 694.26 202.54 695.97 ;
   RECT 23.18 695.97 202.54 697.68 ;
   RECT 23.18 697.68 202.54 699.39 ;
   RECT 23.18 699.39 202.54 701.1 ;
   RECT 23.18 701.1 202.54 702.81 ;
   RECT 23.18 702.81 202.54 704.52 ;
   RECT 23.18 704.52 202.54 706.23 ;
   RECT 23.18 706.23 202.54 707.94 ;
   RECT 23.18 707.94 202.54 709.65 ;
   RECT 23.18 709.65 202.54 711.36 ;
   RECT 23.18 711.36 202.54 713.07 ;
   RECT 23.18 713.07 202.54 714.78 ;
   RECT 23.18 714.78 202.54 716.49 ;
   RECT 23.18 716.49 202.54 718.2 ;
   RECT 23.18 718.2 202.54 719.91 ;
   RECT 23.18 719.91 202.54 721.62 ;
   RECT 23.18 721.62 202.54 723.33 ;
   RECT 23.18 723.33 202.54 725.04 ;
   RECT 23.18 725.04 202.54 726.75 ;
   RECT 23.18 726.75 202.54 728.46 ;
   RECT 23.18 728.46 202.54 730.17 ;
   RECT 23.18 730.17 202.54 731.88 ;
   RECT 23.18 731.88 202.54 733.59 ;
   RECT 23.18 733.59 202.54 735.3 ;
   RECT 23.18 735.3 202.54 737.01 ;
   RECT 23.18 737.01 202.54 738.72 ;
   RECT 23.18 738.72 202.54 740.43 ;
   RECT 23.18 740.43 202.54 742.14 ;
   RECT 23.18 742.14 202.54 743.85 ;
   RECT 23.18 743.85 202.54 745.56 ;
   RECT 23.18 745.56 202.54 747.27 ;
   RECT 23.18 747.27 202.54 748.98 ;
   RECT 23.18 748.98 202.54 750.69 ;
   RECT 23.18 750.69 202.54 752.4 ;
   RECT 23.18 752.4 202.54 754.11 ;
   RECT 23.18 754.11 202.54 755.82 ;
   RECT 23.18 755.82 202.54 757.53 ;
   RECT 23.18 757.53 202.54 759.24 ;
   RECT 23.18 759.24 202.54 760.95 ;
   RECT 23.18 760.95 202.54 762.66 ;
   RECT 23.18 762.66 202.54 764.37 ;
   RECT 23.18 764.37 202.54 766.08 ;
   RECT 23.18 766.08 202.54 767.79 ;
   RECT 23.18 767.79 202.54 769.5 ;
   RECT 23.18 769.5 202.54 771.21 ;
   RECT 23.18 771.21 202.54 772.92 ;
   RECT 23.18 772.92 202.54 774.63 ;
   RECT 23.18 774.63 202.54 776.34 ;
   RECT 23.18 776.34 202.54 778.05 ;
   RECT 23.18 778.05 202.54 779.76 ;
   RECT 23.18 779.76 202.54 781.47 ;
   RECT 23.18 781.47 202.54 783.18 ;
   RECT 23.18 783.18 202.54 784.89 ;
   RECT 23.18 784.89 202.54 786.6 ;
   RECT 23.18 786.6 202.54 788.31 ;
   RECT 23.18 788.31 202.54 790.02 ;
   RECT 23.18 790.02 202.54 791.73 ;
   RECT 23.18 791.73 202.54 793.44 ;
   RECT 23.18 793.44 202.54 795.15 ;
   RECT 23.18 795.15 202.54 796.86 ;
   RECT 23.18 796.86 202.54 798.57 ;
   RECT 23.18 798.57 202.54 800.28 ;
   RECT 23.18 800.28 202.54 801.99 ;
   RECT 23.18 801.99 202.54 803.7 ;
   RECT 23.18 803.7 202.54 805.41 ;
   RECT 23.18 805.41 202.54 807.12 ;
   RECT 23.18 807.12 202.54 808.83 ;
   RECT 23.18 808.83 202.54 810.54 ;
   RECT 23.18 810.54 202.54 812.25 ;
   RECT 23.18 812.25 202.54 813.96 ;
   RECT 23.18 813.96 202.54 815.67 ;
   RECT 23.18 815.67 202.54 817.38 ;
   RECT 23.18 817.38 202.54 819.09 ;
   RECT 23.18 819.09 202.54 820.8 ;
   RECT 23.18 820.8 202.54 822.51 ;
   RECT 23.18 822.51 202.54 824.22 ;
   RECT 23.18 824.22 202.54 825.93 ;
   RECT 23.18 825.93 202.54 827.64 ;
   RECT 23.18 827.64 202.54 829.35 ;
   RECT 23.18 829.35 202.54 831.06 ;
   RECT 23.18 831.06 202.54 832.77 ;
   RECT 23.18 832.77 202.54 834.48 ;
   RECT 23.18 834.48 202.54 836.19 ;
   RECT 23.18 836.19 202.54 837.9 ;
   RECT 23.18 837.9 202.54 839.61 ;
   RECT 23.18 839.61 202.54 841.32 ;
  LAYER via3 ;
   RECT 23.18 0.0 202.54 1.71 ;
   RECT 23.18 1.71 202.54 3.42 ;
   RECT 23.18 3.42 202.54 5.13 ;
   RECT 23.18 5.13 202.54 6.84 ;
   RECT 23.18 6.84 202.54 8.55 ;
   RECT 23.18 8.55 202.54 10.26 ;
   RECT 23.18 10.26 202.54 11.97 ;
   RECT 23.18 11.97 202.54 13.68 ;
   RECT 23.18 13.68 202.54 15.39 ;
   RECT 23.18 15.39 202.54 17.1 ;
   RECT 23.18 17.1 202.54 18.81 ;
   RECT 23.18 18.81 202.54 20.52 ;
   RECT 23.18 20.52 202.54 22.23 ;
   RECT 23.18 22.23 202.54 23.94 ;
   RECT 23.18 23.94 202.54 25.65 ;
   RECT 23.18 25.65 202.54 27.36 ;
   RECT 23.18 27.36 202.54 29.07 ;
   RECT 23.18 29.07 202.54 30.78 ;
   RECT 23.18 30.78 202.54 32.49 ;
   RECT 23.18 32.49 202.54 34.2 ;
   RECT 23.18 34.2 202.54 35.91 ;
   RECT 23.18 35.91 202.54 37.62 ;
   RECT 23.18 37.62 202.54 39.33 ;
   RECT 23.18 39.33 202.54 41.04 ;
   RECT 23.18 41.04 202.54 42.75 ;
   RECT 23.18 42.75 202.54 44.46 ;
   RECT 23.18 44.46 202.54 46.17 ;
   RECT 23.18 46.17 202.54 47.88 ;
   RECT 23.18 47.88 202.54 49.59 ;
   RECT 23.18 49.59 202.54 51.3 ;
   RECT 23.18 51.3 202.54 53.01 ;
   RECT 23.18 53.01 202.54 54.72 ;
   RECT 23.18 54.72 202.54 56.43 ;
   RECT 23.18 56.43 202.54 58.14 ;
   RECT 23.18 58.14 202.54 59.85 ;
   RECT 23.18 59.85 202.54 61.56 ;
   RECT 23.18 61.56 202.54 63.27 ;
   RECT 23.18 63.27 202.54 64.98 ;
   RECT 23.18 64.98 202.54 66.69 ;
   RECT 23.18 66.69 202.54 68.4 ;
   RECT 23.18 68.4 202.54 70.11 ;
   RECT 23.18 70.11 202.54 71.82 ;
   RECT 23.18 71.82 202.54 73.53 ;
   RECT 23.18 73.53 202.54 75.24 ;
   RECT 23.18 75.24 202.54 76.95 ;
   RECT 23.18 76.95 202.54 78.66 ;
   RECT 23.18 78.66 202.54 80.37 ;
   RECT 23.18 80.37 202.54 82.08 ;
   RECT 23.18 82.08 202.54 83.79 ;
   RECT 23.18 83.79 202.54 85.5 ;
   RECT 23.18 85.5 202.54 87.21 ;
   RECT 23.18 87.21 202.54 88.92 ;
   RECT 23.18 88.92 202.54 90.63 ;
   RECT 23.18 90.63 202.54 92.34 ;
   RECT 23.18 92.34 202.54 94.05 ;
   RECT 23.18 94.05 202.54 95.76 ;
   RECT 23.18 95.76 202.54 97.47 ;
   RECT 23.18 97.47 202.54 99.18 ;
   RECT 23.18 99.18 202.54 100.89 ;
   RECT 23.18 100.89 202.54 102.6 ;
   RECT 23.18 102.6 202.54 104.31 ;
   RECT 23.18 104.31 202.54 106.02 ;
   RECT 23.18 106.02 202.54 107.73 ;
   RECT 23.18 107.73 202.54 109.44 ;
   RECT 23.18 109.44 202.54 111.15 ;
   RECT 23.18 111.15 202.54 112.86 ;
   RECT 23.18 112.86 202.54 114.57 ;
   RECT 23.18 114.57 202.54 116.28 ;
   RECT 23.18 116.28 202.54 117.99 ;
   RECT 23.18 117.99 202.54 119.7 ;
   RECT 23.18 119.7 202.54 121.41 ;
   RECT 23.18 121.41 202.54 123.12 ;
   RECT 23.18 123.12 202.54 124.83 ;
   RECT 23.18 124.83 202.54 126.54 ;
   RECT 23.18 126.54 202.54 128.25 ;
   RECT 23.18 128.25 202.54 129.96 ;
   RECT 23.18 129.96 202.54 131.67 ;
   RECT 23.18 131.67 202.54 133.38 ;
   RECT 23.18 133.38 202.54 135.09 ;
   RECT 23.18 135.09 202.54 136.8 ;
   RECT 23.18 136.8 202.54 138.51 ;
   RECT 23.18 138.51 202.54 140.22 ;
   RECT 23.18 140.22 202.54 141.93 ;
   RECT 23.18 141.93 202.54 143.64 ;
   RECT 23.18 143.64 202.54 145.35 ;
   RECT 23.18 145.35 202.54 147.06 ;
   RECT 23.18 147.06 202.54 148.77 ;
   RECT 23.18 148.77 202.54 150.48 ;
   RECT 23.18 150.48 202.54 152.19 ;
   RECT 23.18 152.19 202.54 153.9 ;
   RECT 23.18 153.9 202.54 155.61 ;
   RECT 23.18 155.61 202.54 157.32 ;
   RECT 23.18 157.32 202.54 159.03 ;
   RECT 23.18 159.03 202.54 160.74 ;
   RECT 23.18 160.74 202.54 162.45 ;
   RECT 23.18 162.45 202.54 164.16 ;
   RECT 23.18 164.16 202.54 165.87 ;
   RECT 23.18 165.87 202.54 167.58 ;
   RECT 23.18 167.58 202.54 169.29 ;
   RECT 23.18 169.29 202.54 171.0 ;
   RECT 23.18 171.0 202.54 172.71 ;
   RECT 23.18 172.71 202.54 174.42 ;
   RECT 23.18 174.42 202.54 176.13 ;
   RECT 23.18 176.13 202.54 177.84 ;
   RECT 23.18 177.84 202.54 179.55 ;
   RECT 23.18 179.55 202.54 181.26 ;
   RECT 23.18 181.26 202.54 182.97 ;
   RECT 23.18 182.97 202.54 184.68 ;
   RECT 23.18 184.68 202.54 186.39 ;
   RECT 23.18 186.39 202.54 188.1 ;
   RECT 23.18 188.1 202.54 189.81 ;
   RECT 23.18 189.81 202.54 191.52 ;
   RECT 23.18 191.52 202.54 193.23 ;
   RECT 23.18 193.23 202.54 194.94 ;
   RECT 23.18 194.94 202.54 196.65 ;
   RECT 23.18 196.65 202.54 198.36 ;
   RECT 23.18 198.36 202.54 200.07 ;
   RECT 23.18 200.07 202.54 201.78 ;
   RECT 23.18 201.78 202.54 203.49 ;
   RECT 23.18 203.49 202.54 205.2 ;
   RECT 23.18 205.2 202.54 206.91 ;
   RECT 23.18 206.91 202.54 208.62 ;
   RECT 23.18 208.62 202.54 210.33 ;
   RECT 23.18 210.33 202.54 212.04 ;
   RECT 23.18 212.04 202.54 213.75 ;
   RECT 23.18 213.75 202.54 215.46 ;
   RECT 23.18 215.46 202.54 217.17 ;
   RECT 23.18 217.17 202.54 218.88 ;
   RECT 23.18 218.88 202.54 220.59 ;
   RECT 23.18 220.59 202.54 222.3 ;
   RECT 23.18 222.3 202.54 224.01 ;
   RECT 23.18 224.01 202.54 225.72 ;
   RECT 23.18 225.72 202.54 227.43 ;
   RECT 23.18 227.43 202.54 229.14 ;
   RECT 23.18 229.14 202.54 230.85 ;
   RECT 23.18 230.85 202.54 232.56 ;
   RECT 23.18 232.56 202.54 234.27 ;
   RECT 23.18 234.27 202.54 235.98 ;
   RECT 23.18 235.98 202.54 237.69 ;
   RECT 23.18 237.69 202.54 239.4 ;
   RECT 23.18 239.4 202.54 241.11 ;
   RECT 23.18 241.11 202.54 242.82 ;
   RECT 23.18 242.82 202.54 244.53 ;
   RECT 23.18 244.53 202.54 246.24 ;
   RECT 23.18 246.24 202.54 247.95 ;
   RECT 23.18 247.95 202.54 249.66 ;
   RECT 23.18 249.66 202.54 251.37 ;
   RECT 23.18 251.37 202.54 253.08 ;
   RECT 23.18 253.08 202.54 254.79 ;
   RECT 23.18 254.79 202.54 256.5 ;
   RECT 23.18 256.5 202.54 258.21 ;
   RECT 23.18 258.21 202.54 259.92 ;
   RECT 23.18 259.92 202.54 261.63 ;
   RECT 23.18 261.63 202.54 263.34 ;
   RECT 23.18 263.34 202.54 265.05 ;
   RECT 23.18 265.05 202.54 266.76 ;
   RECT 23.18 266.76 202.54 268.47 ;
   RECT 23.18 268.47 202.54 270.18 ;
   RECT 23.18 270.18 202.54 271.89 ;
   RECT 23.18 271.89 202.54 273.6 ;
   RECT 23.18 273.6 202.54 275.31 ;
   RECT 23.18 275.31 202.54 277.02 ;
   RECT 23.18 277.02 202.54 278.73 ;
   RECT 23.18 278.73 202.54 280.44 ;
   RECT 23.18 280.44 202.54 282.15 ;
   RECT 23.18 282.15 202.54 283.86 ;
   RECT 23.18 283.86 202.54 285.57 ;
   RECT 23.18 285.57 202.54 287.28 ;
   RECT 23.18 287.28 202.54 288.99 ;
   RECT 23.18 288.99 202.54 290.7 ;
   RECT 23.18 290.7 202.54 292.41 ;
   RECT 23.18 292.41 202.54 294.12 ;
   RECT 23.18 294.12 202.54 295.83 ;
   RECT 23.18 295.83 202.54 297.54 ;
   RECT 23.18 297.54 202.54 299.25 ;
   RECT 23.18 299.25 202.54 300.96 ;
   RECT 23.18 300.96 202.54 302.67 ;
   RECT 23.18 302.67 202.54 304.38 ;
   RECT 23.18 304.38 202.54 306.09 ;
   RECT 23.18 306.09 202.54 307.8 ;
   RECT 23.18 307.8 202.54 309.51 ;
   RECT 23.18 309.51 202.54 311.22 ;
   RECT 23.18 311.22 202.54 312.93 ;
   RECT 23.18 312.93 202.54 314.64 ;
   RECT 23.18 314.64 202.54 316.35 ;
   RECT 23.18 316.35 202.54 318.06 ;
   RECT 23.18 318.06 202.54 319.77 ;
   RECT 23.18 319.77 202.54 321.48 ;
   RECT 23.18 321.48 202.54 323.19 ;
   RECT 23.18 323.19 202.54 324.9 ;
   RECT 23.18 324.9 202.54 326.61 ;
   RECT 23.18 326.61 202.54 328.32 ;
   RECT 23.18 328.32 202.54 330.03 ;
   RECT 23.18 330.03 202.54 331.74 ;
   RECT 23.18 331.74 202.54 333.45 ;
   RECT 23.18 333.45 202.54 335.16 ;
   RECT 23.18 335.16 202.54 336.87 ;
   RECT 23.18 336.87 202.54 338.58 ;
   RECT 23.18 338.58 202.54 340.29 ;
   RECT 23.18 340.29 202.54 342.0 ;
   RECT 23.18 342.0 202.54 343.71 ;
   RECT 23.18 343.71 202.54 345.42 ;
   RECT 23.18 345.42 202.54 347.13 ;
   RECT 23.18 347.13 202.54 348.84 ;
   RECT 23.18 348.84 202.54 350.55 ;
   RECT 23.18 350.55 202.54 352.26 ;
   RECT 23.18 352.26 202.54 353.97 ;
   RECT 23.18 353.97 202.54 355.68 ;
   RECT 23.18 355.68 202.54 357.39 ;
   RECT 23.18 357.39 202.54 359.1 ;
   RECT 23.18 359.1 202.54 360.81 ;
   RECT 23.18 360.81 202.54 362.52 ;
   RECT 23.18 362.52 202.54 364.23 ;
   RECT 23.18 364.23 202.54 365.94 ;
   RECT 23.18 365.94 202.54 367.65 ;
   RECT 23.18 367.65 202.54 369.36 ;
   RECT 23.18 369.36 202.54 371.07 ;
   RECT 23.18 371.07 202.54 372.78 ;
   RECT 23.18 372.78 202.54 374.49 ;
   RECT 23.18 374.49 202.54 376.2 ;
   RECT 23.18 376.2 202.54 377.91 ;
   RECT 23.18 377.91 202.54 379.62 ;
   RECT 23.18 379.62 202.54 381.33 ;
   RECT 23.18 381.33 202.54 383.04 ;
   RECT 23.18 383.04 202.54 384.75 ;
   RECT 23.18 384.75 202.54 386.46 ;
   RECT 23.18 386.46 202.54 388.17 ;
   RECT 23.18 388.17 202.54 389.88 ;
   RECT 23.18 389.88 202.54 391.59 ;
   RECT 23.18 391.59 202.54 393.3 ;
   RECT 23.18 393.3 202.54 395.01 ;
   RECT 23.18 395.01 202.54 396.72 ;
   RECT 23.18 396.72 202.54 398.43 ;
   RECT 23.18 398.43 202.54 400.14 ;
   RECT 23.18 400.14 202.54 401.85 ;
   RECT 0.0 401.85 202.54 403.56 ;
   RECT 0.0 403.56 202.54 405.27 ;
   RECT 0.0 405.27 202.54 406.98 ;
   RECT 0.0 406.98 202.54 408.69 ;
   RECT 0.0 408.69 202.54 410.4 ;
   RECT 0.0 410.4 202.54 412.11 ;
   RECT 0.0 412.11 202.54 413.82 ;
   RECT 0.0 413.82 202.54 415.53 ;
   RECT 0.0 415.53 202.54 417.24 ;
   RECT 0.0 417.24 202.54 418.95 ;
   RECT 0.0 418.95 202.54 420.66 ;
   RECT 0.0 420.66 202.54 422.37 ;
   RECT 0.0 422.37 202.54 424.08 ;
   RECT 0.0 424.08 202.54 425.79 ;
   RECT 0.0 425.79 202.54 427.5 ;
   RECT 0.0 427.5 202.54 429.21 ;
   RECT 0.0 429.21 202.54 430.92 ;
   RECT 23.18 430.92 202.54 432.63 ;
   RECT 23.18 432.63 202.54 434.34 ;
   RECT 23.18 434.34 202.54 436.05 ;
   RECT 23.18 436.05 202.54 437.76 ;
   RECT 23.18 437.76 202.54 439.47 ;
   RECT 23.18 439.47 202.54 441.18 ;
   RECT 23.18 441.18 202.54 442.89 ;
   RECT 23.18 442.89 202.54 444.6 ;
   RECT 23.18 444.6 202.54 446.31 ;
   RECT 23.18 446.31 202.54 448.02 ;
   RECT 23.18 448.02 202.54 449.73 ;
   RECT 23.18 449.73 202.54 451.44 ;
   RECT 23.18 451.44 202.54 453.15 ;
   RECT 23.18 453.15 202.54 454.86 ;
   RECT 23.18 454.86 202.54 456.57 ;
   RECT 23.18 456.57 202.54 458.28 ;
   RECT 23.18 458.28 202.54 459.99 ;
   RECT 23.18 459.99 202.54 461.7 ;
   RECT 23.18 461.7 202.54 463.41 ;
   RECT 23.18 463.41 202.54 465.12 ;
   RECT 23.18 465.12 202.54 466.83 ;
   RECT 23.18 466.83 202.54 468.54 ;
   RECT 23.18 468.54 202.54 470.25 ;
   RECT 23.18 470.25 202.54 471.96 ;
   RECT 23.18 471.96 202.54 473.67 ;
   RECT 23.18 473.67 202.54 475.38 ;
   RECT 23.18 475.38 202.54 477.09 ;
   RECT 23.18 477.09 202.54 478.8 ;
   RECT 23.18 478.8 202.54 480.51 ;
   RECT 23.18 480.51 202.54 482.22 ;
   RECT 23.18 482.22 202.54 483.93 ;
   RECT 23.18 483.93 202.54 485.64 ;
   RECT 23.18 485.64 202.54 487.35 ;
   RECT 23.18 487.35 202.54 489.06 ;
   RECT 23.18 489.06 202.54 490.77 ;
   RECT 23.18 490.77 202.54 492.48 ;
   RECT 23.18 492.48 202.54 494.19 ;
   RECT 23.18 494.19 202.54 495.9 ;
   RECT 23.18 495.9 202.54 497.61 ;
   RECT 23.18 497.61 202.54 499.32 ;
   RECT 23.18 499.32 202.54 501.03 ;
   RECT 23.18 501.03 202.54 502.74 ;
   RECT 23.18 502.74 202.54 504.45 ;
   RECT 23.18 504.45 202.54 506.16 ;
   RECT 23.18 506.16 202.54 507.87 ;
   RECT 23.18 507.87 202.54 509.58 ;
   RECT 23.18 509.58 202.54 511.29 ;
   RECT 23.18 511.29 202.54 513.0 ;
   RECT 23.18 513.0 202.54 514.71 ;
   RECT 23.18 514.71 202.54 516.42 ;
   RECT 23.18 516.42 202.54 518.13 ;
   RECT 23.18 518.13 202.54 519.84 ;
   RECT 23.18 519.84 202.54 521.55 ;
   RECT 23.18 521.55 202.54 523.26 ;
   RECT 23.18 523.26 202.54 524.97 ;
   RECT 23.18 524.97 202.54 526.68 ;
   RECT 23.18 526.68 202.54 528.39 ;
   RECT 23.18 528.39 202.54 530.1 ;
   RECT 23.18 530.1 202.54 531.81 ;
   RECT 23.18 531.81 202.54 533.52 ;
   RECT 23.18 533.52 202.54 535.23 ;
   RECT 23.18 535.23 202.54 536.94 ;
   RECT 23.18 536.94 202.54 538.65 ;
   RECT 23.18 538.65 202.54 540.36 ;
   RECT 23.18 540.36 202.54 542.07 ;
   RECT 23.18 542.07 202.54 543.78 ;
   RECT 23.18 543.78 202.54 545.49 ;
   RECT 23.18 545.49 202.54 547.2 ;
   RECT 23.18 547.2 202.54 548.91 ;
   RECT 23.18 548.91 202.54 550.62 ;
   RECT 23.18 550.62 202.54 552.33 ;
   RECT 23.18 552.33 202.54 554.04 ;
   RECT 23.18 554.04 202.54 555.75 ;
   RECT 23.18 555.75 202.54 557.46 ;
   RECT 23.18 557.46 202.54 559.17 ;
   RECT 23.18 559.17 202.54 560.88 ;
   RECT 23.18 560.88 202.54 562.59 ;
   RECT 23.18 562.59 202.54 564.3 ;
   RECT 23.18 564.3 202.54 566.01 ;
   RECT 23.18 566.01 202.54 567.72 ;
   RECT 23.18 567.72 202.54 569.43 ;
   RECT 23.18 569.43 202.54 571.14 ;
   RECT 23.18 571.14 202.54 572.85 ;
   RECT 23.18 572.85 202.54 574.56 ;
   RECT 23.18 574.56 202.54 576.27 ;
   RECT 23.18 576.27 202.54 577.98 ;
   RECT 23.18 577.98 202.54 579.69 ;
   RECT 23.18 579.69 202.54 581.4 ;
   RECT 23.18 581.4 202.54 583.11 ;
   RECT 23.18 583.11 202.54 584.82 ;
   RECT 23.18 584.82 202.54 586.53 ;
   RECT 23.18 586.53 202.54 588.24 ;
   RECT 23.18 588.24 202.54 589.95 ;
   RECT 23.18 589.95 202.54 591.66 ;
   RECT 23.18 591.66 202.54 593.37 ;
   RECT 23.18 593.37 202.54 595.08 ;
   RECT 23.18 595.08 202.54 596.79 ;
   RECT 23.18 596.79 202.54 598.5 ;
   RECT 23.18 598.5 202.54 600.21 ;
   RECT 23.18 600.21 202.54 601.92 ;
   RECT 23.18 601.92 202.54 603.63 ;
   RECT 23.18 603.63 202.54 605.34 ;
   RECT 23.18 605.34 202.54 607.05 ;
   RECT 23.18 607.05 202.54 608.76 ;
   RECT 23.18 608.76 202.54 610.47 ;
   RECT 23.18 610.47 202.54 612.18 ;
   RECT 23.18 612.18 202.54 613.89 ;
   RECT 23.18 613.89 202.54 615.6 ;
   RECT 23.18 615.6 202.54 617.31 ;
   RECT 23.18 617.31 202.54 619.02 ;
   RECT 23.18 619.02 202.54 620.73 ;
   RECT 23.18 620.73 202.54 622.44 ;
   RECT 23.18 622.44 202.54 624.15 ;
   RECT 23.18 624.15 202.54 625.86 ;
   RECT 23.18 625.86 202.54 627.57 ;
   RECT 23.18 627.57 202.54 629.28 ;
   RECT 23.18 629.28 202.54 630.99 ;
   RECT 23.18 630.99 202.54 632.7 ;
   RECT 23.18 632.7 202.54 634.41 ;
   RECT 23.18 634.41 202.54 636.12 ;
   RECT 23.18 636.12 202.54 637.83 ;
   RECT 23.18 637.83 202.54 639.54 ;
   RECT 23.18 639.54 202.54 641.25 ;
   RECT 23.18 641.25 202.54 642.96 ;
   RECT 23.18 642.96 202.54 644.67 ;
   RECT 23.18 644.67 202.54 646.38 ;
   RECT 23.18 646.38 202.54 648.09 ;
   RECT 23.18 648.09 202.54 649.8 ;
   RECT 23.18 649.8 202.54 651.51 ;
   RECT 23.18 651.51 202.54 653.22 ;
   RECT 23.18 653.22 202.54 654.93 ;
   RECT 23.18 654.93 202.54 656.64 ;
   RECT 23.18 656.64 202.54 658.35 ;
   RECT 23.18 658.35 202.54 660.06 ;
   RECT 23.18 660.06 202.54 661.77 ;
   RECT 23.18 661.77 202.54 663.48 ;
   RECT 23.18 663.48 202.54 665.19 ;
   RECT 23.18 665.19 202.54 666.9 ;
   RECT 23.18 666.9 202.54 668.61 ;
   RECT 23.18 668.61 202.54 670.32 ;
   RECT 23.18 670.32 202.54 672.03 ;
   RECT 23.18 672.03 202.54 673.74 ;
   RECT 23.18 673.74 202.54 675.45 ;
   RECT 23.18 675.45 202.54 677.16 ;
   RECT 23.18 677.16 202.54 678.87 ;
   RECT 23.18 678.87 202.54 680.58 ;
   RECT 23.18 680.58 202.54 682.29 ;
   RECT 23.18 682.29 202.54 684.0 ;
   RECT 23.18 684.0 202.54 685.71 ;
   RECT 23.18 685.71 202.54 687.42 ;
   RECT 23.18 687.42 202.54 689.13 ;
   RECT 23.18 689.13 202.54 690.84 ;
   RECT 23.18 690.84 202.54 692.55 ;
   RECT 23.18 692.55 202.54 694.26 ;
   RECT 23.18 694.26 202.54 695.97 ;
   RECT 23.18 695.97 202.54 697.68 ;
   RECT 23.18 697.68 202.54 699.39 ;
   RECT 23.18 699.39 202.54 701.1 ;
   RECT 23.18 701.1 202.54 702.81 ;
   RECT 23.18 702.81 202.54 704.52 ;
   RECT 23.18 704.52 202.54 706.23 ;
   RECT 23.18 706.23 202.54 707.94 ;
   RECT 23.18 707.94 202.54 709.65 ;
   RECT 23.18 709.65 202.54 711.36 ;
   RECT 23.18 711.36 202.54 713.07 ;
   RECT 23.18 713.07 202.54 714.78 ;
   RECT 23.18 714.78 202.54 716.49 ;
   RECT 23.18 716.49 202.54 718.2 ;
   RECT 23.18 718.2 202.54 719.91 ;
   RECT 23.18 719.91 202.54 721.62 ;
   RECT 23.18 721.62 202.54 723.33 ;
   RECT 23.18 723.33 202.54 725.04 ;
   RECT 23.18 725.04 202.54 726.75 ;
   RECT 23.18 726.75 202.54 728.46 ;
   RECT 23.18 728.46 202.54 730.17 ;
   RECT 23.18 730.17 202.54 731.88 ;
   RECT 23.18 731.88 202.54 733.59 ;
   RECT 23.18 733.59 202.54 735.3 ;
   RECT 23.18 735.3 202.54 737.01 ;
   RECT 23.18 737.01 202.54 738.72 ;
   RECT 23.18 738.72 202.54 740.43 ;
   RECT 23.18 740.43 202.54 742.14 ;
   RECT 23.18 742.14 202.54 743.85 ;
   RECT 23.18 743.85 202.54 745.56 ;
   RECT 23.18 745.56 202.54 747.27 ;
   RECT 23.18 747.27 202.54 748.98 ;
   RECT 23.18 748.98 202.54 750.69 ;
   RECT 23.18 750.69 202.54 752.4 ;
   RECT 23.18 752.4 202.54 754.11 ;
   RECT 23.18 754.11 202.54 755.82 ;
   RECT 23.18 755.82 202.54 757.53 ;
   RECT 23.18 757.53 202.54 759.24 ;
   RECT 23.18 759.24 202.54 760.95 ;
   RECT 23.18 760.95 202.54 762.66 ;
   RECT 23.18 762.66 202.54 764.37 ;
   RECT 23.18 764.37 202.54 766.08 ;
   RECT 23.18 766.08 202.54 767.79 ;
   RECT 23.18 767.79 202.54 769.5 ;
   RECT 23.18 769.5 202.54 771.21 ;
   RECT 23.18 771.21 202.54 772.92 ;
   RECT 23.18 772.92 202.54 774.63 ;
   RECT 23.18 774.63 202.54 776.34 ;
   RECT 23.18 776.34 202.54 778.05 ;
   RECT 23.18 778.05 202.54 779.76 ;
   RECT 23.18 779.76 202.54 781.47 ;
   RECT 23.18 781.47 202.54 783.18 ;
   RECT 23.18 783.18 202.54 784.89 ;
   RECT 23.18 784.89 202.54 786.6 ;
   RECT 23.18 786.6 202.54 788.31 ;
   RECT 23.18 788.31 202.54 790.02 ;
   RECT 23.18 790.02 202.54 791.73 ;
   RECT 23.18 791.73 202.54 793.44 ;
   RECT 23.18 793.44 202.54 795.15 ;
   RECT 23.18 795.15 202.54 796.86 ;
   RECT 23.18 796.86 202.54 798.57 ;
   RECT 23.18 798.57 202.54 800.28 ;
   RECT 23.18 800.28 202.54 801.99 ;
   RECT 23.18 801.99 202.54 803.7 ;
   RECT 23.18 803.7 202.54 805.41 ;
   RECT 23.18 805.41 202.54 807.12 ;
   RECT 23.18 807.12 202.54 808.83 ;
   RECT 23.18 808.83 202.54 810.54 ;
   RECT 23.18 810.54 202.54 812.25 ;
   RECT 23.18 812.25 202.54 813.96 ;
   RECT 23.18 813.96 202.54 815.67 ;
   RECT 23.18 815.67 202.54 817.38 ;
   RECT 23.18 817.38 202.54 819.09 ;
   RECT 23.18 819.09 202.54 820.8 ;
   RECT 23.18 820.8 202.54 822.51 ;
   RECT 23.18 822.51 202.54 824.22 ;
   RECT 23.18 824.22 202.54 825.93 ;
   RECT 23.18 825.93 202.54 827.64 ;
   RECT 23.18 827.64 202.54 829.35 ;
   RECT 23.18 829.35 202.54 831.06 ;
   RECT 23.18 831.06 202.54 832.77 ;
   RECT 23.18 832.77 202.54 834.48 ;
   RECT 23.18 834.48 202.54 836.19 ;
   RECT 23.18 836.19 202.54 837.9 ;
   RECT 23.18 837.9 202.54 839.61 ;
   RECT 23.18 839.61 202.54 841.32 ;
  LAYER metal4 ;
   RECT 23.18 0.0 202.54 1.71 ;
   RECT 23.18 1.71 202.54 3.42 ;
   RECT 23.18 3.42 202.54 5.13 ;
   RECT 23.18 5.13 202.54 6.84 ;
   RECT 23.18 6.84 202.54 8.55 ;
   RECT 23.18 8.55 202.54 10.26 ;
   RECT 23.18 10.26 202.54 11.97 ;
   RECT 23.18 11.97 202.54 13.68 ;
   RECT 23.18 13.68 202.54 15.39 ;
   RECT 23.18 15.39 202.54 17.1 ;
   RECT 23.18 17.1 202.54 18.81 ;
   RECT 23.18 18.81 202.54 20.52 ;
   RECT 23.18 20.52 202.54 22.23 ;
   RECT 23.18 22.23 202.54 23.94 ;
   RECT 23.18 23.94 202.54 25.65 ;
   RECT 23.18 25.65 202.54 27.36 ;
   RECT 23.18 27.36 202.54 29.07 ;
   RECT 23.18 29.07 202.54 30.78 ;
   RECT 23.18 30.78 202.54 32.49 ;
   RECT 23.18 32.49 202.54 34.2 ;
   RECT 23.18 34.2 202.54 35.91 ;
   RECT 23.18 35.91 202.54 37.62 ;
   RECT 23.18 37.62 202.54 39.33 ;
   RECT 23.18 39.33 202.54 41.04 ;
   RECT 23.18 41.04 202.54 42.75 ;
   RECT 23.18 42.75 202.54 44.46 ;
   RECT 23.18 44.46 202.54 46.17 ;
   RECT 23.18 46.17 202.54 47.88 ;
   RECT 23.18 47.88 202.54 49.59 ;
   RECT 23.18 49.59 202.54 51.3 ;
   RECT 23.18 51.3 202.54 53.01 ;
   RECT 23.18 53.01 202.54 54.72 ;
   RECT 23.18 54.72 202.54 56.43 ;
   RECT 23.18 56.43 202.54 58.14 ;
   RECT 23.18 58.14 202.54 59.85 ;
   RECT 23.18 59.85 202.54 61.56 ;
   RECT 23.18 61.56 202.54 63.27 ;
   RECT 23.18 63.27 202.54 64.98 ;
   RECT 23.18 64.98 202.54 66.69 ;
   RECT 23.18 66.69 202.54 68.4 ;
   RECT 23.18 68.4 202.54 70.11 ;
   RECT 23.18 70.11 202.54 71.82 ;
   RECT 23.18 71.82 202.54 73.53 ;
   RECT 23.18 73.53 202.54 75.24 ;
   RECT 23.18 75.24 202.54 76.95 ;
   RECT 23.18 76.95 202.54 78.66 ;
   RECT 23.18 78.66 202.54 80.37 ;
   RECT 23.18 80.37 202.54 82.08 ;
   RECT 23.18 82.08 202.54 83.79 ;
   RECT 23.18 83.79 202.54 85.5 ;
   RECT 23.18 85.5 202.54 87.21 ;
   RECT 23.18 87.21 202.54 88.92 ;
   RECT 23.18 88.92 202.54 90.63 ;
   RECT 23.18 90.63 202.54 92.34 ;
   RECT 23.18 92.34 202.54 94.05 ;
   RECT 23.18 94.05 202.54 95.76 ;
   RECT 23.18 95.76 202.54 97.47 ;
   RECT 23.18 97.47 202.54 99.18 ;
   RECT 23.18 99.18 202.54 100.89 ;
   RECT 23.18 100.89 202.54 102.6 ;
   RECT 23.18 102.6 202.54 104.31 ;
   RECT 23.18 104.31 202.54 106.02 ;
   RECT 23.18 106.02 202.54 107.73 ;
   RECT 23.18 107.73 202.54 109.44 ;
   RECT 23.18 109.44 202.54 111.15 ;
   RECT 23.18 111.15 202.54 112.86 ;
   RECT 23.18 112.86 202.54 114.57 ;
   RECT 23.18 114.57 202.54 116.28 ;
   RECT 23.18 116.28 202.54 117.99 ;
   RECT 23.18 117.99 202.54 119.7 ;
   RECT 23.18 119.7 202.54 121.41 ;
   RECT 23.18 121.41 202.54 123.12 ;
   RECT 23.18 123.12 202.54 124.83 ;
   RECT 23.18 124.83 202.54 126.54 ;
   RECT 23.18 126.54 202.54 128.25 ;
   RECT 23.18 128.25 202.54 129.96 ;
   RECT 23.18 129.96 202.54 131.67 ;
   RECT 23.18 131.67 202.54 133.38 ;
   RECT 23.18 133.38 202.54 135.09 ;
   RECT 23.18 135.09 202.54 136.8 ;
   RECT 23.18 136.8 202.54 138.51 ;
   RECT 23.18 138.51 202.54 140.22 ;
   RECT 23.18 140.22 202.54 141.93 ;
   RECT 23.18 141.93 202.54 143.64 ;
   RECT 23.18 143.64 202.54 145.35 ;
   RECT 23.18 145.35 202.54 147.06 ;
   RECT 23.18 147.06 202.54 148.77 ;
   RECT 23.18 148.77 202.54 150.48 ;
   RECT 23.18 150.48 202.54 152.19 ;
   RECT 23.18 152.19 202.54 153.9 ;
   RECT 23.18 153.9 202.54 155.61 ;
   RECT 23.18 155.61 202.54 157.32 ;
   RECT 23.18 157.32 202.54 159.03 ;
   RECT 23.18 159.03 202.54 160.74 ;
   RECT 23.18 160.74 202.54 162.45 ;
   RECT 23.18 162.45 202.54 164.16 ;
   RECT 23.18 164.16 202.54 165.87 ;
   RECT 23.18 165.87 202.54 167.58 ;
   RECT 23.18 167.58 202.54 169.29 ;
   RECT 23.18 169.29 202.54 171.0 ;
   RECT 23.18 171.0 202.54 172.71 ;
   RECT 23.18 172.71 202.54 174.42 ;
   RECT 23.18 174.42 202.54 176.13 ;
   RECT 23.18 176.13 202.54 177.84 ;
   RECT 23.18 177.84 202.54 179.55 ;
   RECT 23.18 179.55 202.54 181.26 ;
   RECT 23.18 181.26 202.54 182.97 ;
   RECT 23.18 182.97 202.54 184.68 ;
   RECT 23.18 184.68 202.54 186.39 ;
   RECT 23.18 186.39 202.54 188.1 ;
   RECT 23.18 188.1 202.54 189.81 ;
   RECT 23.18 189.81 202.54 191.52 ;
   RECT 23.18 191.52 202.54 193.23 ;
   RECT 23.18 193.23 202.54 194.94 ;
   RECT 23.18 194.94 202.54 196.65 ;
   RECT 23.18 196.65 202.54 198.36 ;
   RECT 23.18 198.36 202.54 200.07 ;
   RECT 23.18 200.07 202.54 201.78 ;
   RECT 23.18 201.78 202.54 203.49 ;
   RECT 23.18 203.49 202.54 205.2 ;
   RECT 23.18 205.2 202.54 206.91 ;
   RECT 23.18 206.91 202.54 208.62 ;
   RECT 23.18 208.62 202.54 210.33 ;
   RECT 23.18 210.33 202.54 212.04 ;
   RECT 23.18 212.04 202.54 213.75 ;
   RECT 23.18 213.75 202.54 215.46 ;
   RECT 23.18 215.46 202.54 217.17 ;
   RECT 23.18 217.17 202.54 218.88 ;
   RECT 23.18 218.88 202.54 220.59 ;
   RECT 23.18 220.59 202.54 222.3 ;
   RECT 23.18 222.3 202.54 224.01 ;
   RECT 23.18 224.01 202.54 225.72 ;
   RECT 23.18 225.72 202.54 227.43 ;
   RECT 23.18 227.43 202.54 229.14 ;
   RECT 23.18 229.14 202.54 230.85 ;
   RECT 23.18 230.85 202.54 232.56 ;
   RECT 23.18 232.56 202.54 234.27 ;
   RECT 23.18 234.27 202.54 235.98 ;
   RECT 23.18 235.98 202.54 237.69 ;
   RECT 23.18 237.69 202.54 239.4 ;
   RECT 23.18 239.4 202.54 241.11 ;
   RECT 23.18 241.11 202.54 242.82 ;
   RECT 23.18 242.82 202.54 244.53 ;
   RECT 23.18 244.53 202.54 246.24 ;
   RECT 23.18 246.24 202.54 247.95 ;
   RECT 23.18 247.95 202.54 249.66 ;
   RECT 23.18 249.66 202.54 251.37 ;
   RECT 23.18 251.37 202.54 253.08 ;
   RECT 23.18 253.08 202.54 254.79 ;
   RECT 23.18 254.79 202.54 256.5 ;
   RECT 23.18 256.5 202.54 258.21 ;
   RECT 23.18 258.21 202.54 259.92 ;
   RECT 23.18 259.92 202.54 261.63 ;
   RECT 23.18 261.63 202.54 263.34 ;
   RECT 23.18 263.34 202.54 265.05 ;
   RECT 23.18 265.05 202.54 266.76 ;
   RECT 23.18 266.76 202.54 268.47 ;
   RECT 23.18 268.47 202.54 270.18 ;
   RECT 23.18 270.18 202.54 271.89 ;
   RECT 23.18 271.89 202.54 273.6 ;
   RECT 23.18 273.6 202.54 275.31 ;
   RECT 23.18 275.31 202.54 277.02 ;
   RECT 23.18 277.02 202.54 278.73 ;
   RECT 23.18 278.73 202.54 280.44 ;
   RECT 23.18 280.44 202.54 282.15 ;
   RECT 23.18 282.15 202.54 283.86 ;
   RECT 23.18 283.86 202.54 285.57 ;
   RECT 23.18 285.57 202.54 287.28 ;
   RECT 23.18 287.28 202.54 288.99 ;
   RECT 23.18 288.99 202.54 290.7 ;
   RECT 23.18 290.7 202.54 292.41 ;
   RECT 23.18 292.41 202.54 294.12 ;
   RECT 23.18 294.12 202.54 295.83 ;
   RECT 23.18 295.83 202.54 297.54 ;
   RECT 23.18 297.54 202.54 299.25 ;
   RECT 23.18 299.25 202.54 300.96 ;
   RECT 23.18 300.96 202.54 302.67 ;
   RECT 23.18 302.67 202.54 304.38 ;
   RECT 23.18 304.38 202.54 306.09 ;
   RECT 23.18 306.09 202.54 307.8 ;
   RECT 23.18 307.8 202.54 309.51 ;
   RECT 23.18 309.51 202.54 311.22 ;
   RECT 23.18 311.22 202.54 312.93 ;
   RECT 23.18 312.93 202.54 314.64 ;
   RECT 23.18 314.64 202.54 316.35 ;
   RECT 23.18 316.35 202.54 318.06 ;
   RECT 23.18 318.06 202.54 319.77 ;
   RECT 23.18 319.77 202.54 321.48 ;
   RECT 23.18 321.48 202.54 323.19 ;
   RECT 23.18 323.19 202.54 324.9 ;
   RECT 23.18 324.9 202.54 326.61 ;
   RECT 23.18 326.61 202.54 328.32 ;
   RECT 23.18 328.32 202.54 330.03 ;
   RECT 23.18 330.03 202.54 331.74 ;
   RECT 23.18 331.74 202.54 333.45 ;
   RECT 23.18 333.45 202.54 335.16 ;
   RECT 23.18 335.16 202.54 336.87 ;
   RECT 23.18 336.87 202.54 338.58 ;
   RECT 23.18 338.58 202.54 340.29 ;
   RECT 23.18 340.29 202.54 342.0 ;
   RECT 23.18 342.0 202.54 343.71 ;
   RECT 23.18 343.71 202.54 345.42 ;
   RECT 23.18 345.42 202.54 347.13 ;
   RECT 23.18 347.13 202.54 348.84 ;
   RECT 23.18 348.84 202.54 350.55 ;
   RECT 23.18 350.55 202.54 352.26 ;
   RECT 23.18 352.26 202.54 353.97 ;
   RECT 23.18 353.97 202.54 355.68 ;
   RECT 23.18 355.68 202.54 357.39 ;
   RECT 23.18 357.39 202.54 359.1 ;
   RECT 23.18 359.1 202.54 360.81 ;
   RECT 23.18 360.81 202.54 362.52 ;
   RECT 23.18 362.52 202.54 364.23 ;
   RECT 23.18 364.23 202.54 365.94 ;
   RECT 23.18 365.94 202.54 367.65 ;
   RECT 23.18 367.65 202.54 369.36 ;
   RECT 23.18 369.36 202.54 371.07 ;
   RECT 23.18 371.07 202.54 372.78 ;
   RECT 23.18 372.78 202.54 374.49 ;
   RECT 23.18 374.49 202.54 376.2 ;
   RECT 23.18 376.2 202.54 377.91 ;
   RECT 23.18 377.91 202.54 379.62 ;
   RECT 23.18 379.62 202.54 381.33 ;
   RECT 23.18 381.33 202.54 383.04 ;
   RECT 23.18 383.04 202.54 384.75 ;
   RECT 23.18 384.75 202.54 386.46 ;
   RECT 23.18 386.46 202.54 388.17 ;
   RECT 23.18 388.17 202.54 389.88 ;
   RECT 23.18 389.88 202.54 391.59 ;
   RECT 23.18 391.59 202.54 393.3 ;
   RECT 23.18 393.3 202.54 395.01 ;
   RECT 23.18 395.01 202.54 396.72 ;
   RECT 23.18 396.72 202.54 398.43 ;
   RECT 23.18 398.43 202.54 400.14 ;
   RECT 23.18 400.14 202.54 401.85 ;
   RECT 0.0 401.85 202.54 403.56 ;
   RECT 0.0 403.56 202.54 405.27 ;
   RECT 0.0 405.27 202.54 406.98 ;
   RECT 0.0 406.98 202.54 408.69 ;
   RECT 0.0 408.69 202.54 410.4 ;
   RECT 0.0 410.4 202.54 412.11 ;
   RECT 0.0 412.11 202.54 413.82 ;
   RECT 0.0 413.82 202.54 415.53 ;
   RECT 0.0 415.53 202.54 417.24 ;
   RECT 0.0 417.24 202.54 418.95 ;
   RECT 0.0 418.95 202.54 420.66 ;
   RECT 0.0 420.66 202.54 422.37 ;
   RECT 0.0 422.37 202.54 424.08 ;
   RECT 0.0 424.08 202.54 425.79 ;
   RECT 0.0 425.79 202.54 427.5 ;
   RECT 0.0 427.5 202.54 429.21 ;
   RECT 0.0 429.21 202.54 430.92 ;
   RECT 23.18 430.92 202.54 432.63 ;
   RECT 23.18 432.63 202.54 434.34 ;
   RECT 23.18 434.34 202.54 436.05 ;
   RECT 23.18 436.05 202.54 437.76 ;
   RECT 23.18 437.76 202.54 439.47 ;
   RECT 23.18 439.47 202.54 441.18 ;
   RECT 23.18 441.18 202.54 442.89 ;
   RECT 23.18 442.89 202.54 444.6 ;
   RECT 23.18 444.6 202.54 446.31 ;
   RECT 23.18 446.31 202.54 448.02 ;
   RECT 23.18 448.02 202.54 449.73 ;
   RECT 23.18 449.73 202.54 451.44 ;
   RECT 23.18 451.44 202.54 453.15 ;
   RECT 23.18 453.15 202.54 454.86 ;
   RECT 23.18 454.86 202.54 456.57 ;
   RECT 23.18 456.57 202.54 458.28 ;
   RECT 23.18 458.28 202.54 459.99 ;
   RECT 23.18 459.99 202.54 461.7 ;
   RECT 23.18 461.7 202.54 463.41 ;
   RECT 23.18 463.41 202.54 465.12 ;
   RECT 23.18 465.12 202.54 466.83 ;
   RECT 23.18 466.83 202.54 468.54 ;
   RECT 23.18 468.54 202.54 470.25 ;
   RECT 23.18 470.25 202.54 471.96 ;
   RECT 23.18 471.96 202.54 473.67 ;
   RECT 23.18 473.67 202.54 475.38 ;
   RECT 23.18 475.38 202.54 477.09 ;
   RECT 23.18 477.09 202.54 478.8 ;
   RECT 23.18 478.8 202.54 480.51 ;
   RECT 23.18 480.51 202.54 482.22 ;
   RECT 23.18 482.22 202.54 483.93 ;
   RECT 23.18 483.93 202.54 485.64 ;
   RECT 23.18 485.64 202.54 487.35 ;
   RECT 23.18 487.35 202.54 489.06 ;
   RECT 23.18 489.06 202.54 490.77 ;
   RECT 23.18 490.77 202.54 492.48 ;
   RECT 23.18 492.48 202.54 494.19 ;
   RECT 23.18 494.19 202.54 495.9 ;
   RECT 23.18 495.9 202.54 497.61 ;
   RECT 23.18 497.61 202.54 499.32 ;
   RECT 23.18 499.32 202.54 501.03 ;
   RECT 23.18 501.03 202.54 502.74 ;
   RECT 23.18 502.74 202.54 504.45 ;
   RECT 23.18 504.45 202.54 506.16 ;
   RECT 23.18 506.16 202.54 507.87 ;
   RECT 23.18 507.87 202.54 509.58 ;
   RECT 23.18 509.58 202.54 511.29 ;
   RECT 23.18 511.29 202.54 513.0 ;
   RECT 23.18 513.0 202.54 514.71 ;
   RECT 23.18 514.71 202.54 516.42 ;
   RECT 23.18 516.42 202.54 518.13 ;
   RECT 23.18 518.13 202.54 519.84 ;
   RECT 23.18 519.84 202.54 521.55 ;
   RECT 23.18 521.55 202.54 523.26 ;
   RECT 23.18 523.26 202.54 524.97 ;
   RECT 23.18 524.97 202.54 526.68 ;
   RECT 23.18 526.68 202.54 528.39 ;
   RECT 23.18 528.39 202.54 530.1 ;
   RECT 23.18 530.1 202.54 531.81 ;
   RECT 23.18 531.81 202.54 533.52 ;
   RECT 23.18 533.52 202.54 535.23 ;
   RECT 23.18 535.23 202.54 536.94 ;
   RECT 23.18 536.94 202.54 538.65 ;
   RECT 23.18 538.65 202.54 540.36 ;
   RECT 23.18 540.36 202.54 542.07 ;
   RECT 23.18 542.07 202.54 543.78 ;
   RECT 23.18 543.78 202.54 545.49 ;
   RECT 23.18 545.49 202.54 547.2 ;
   RECT 23.18 547.2 202.54 548.91 ;
   RECT 23.18 548.91 202.54 550.62 ;
   RECT 23.18 550.62 202.54 552.33 ;
   RECT 23.18 552.33 202.54 554.04 ;
   RECT 23.18 554.04 202.54 555.75 ;
   RECT 23.18 555.75 202.54 557.46 ;
   RECT 23.18 557.46 202.54 559.17 ;
   RECT 23.18 559.17 202.54 560.88 ;
   RECT 23.18 560.88 202.54 562.59 ;
   RECT 23.18 562.59 202.54 564.3 ;
   RECT 23.18 564.3 202.54 566.01 ;
   RECT 23.18 566.01 202.54 567.72 ;
   RECT 23.18 567.72 202.54 569.43 ;
   RECT 23.18 569.43 202.54 571.14 ;
   RECT 23.18 571.14 202.54 572.85 ;
   RECT 23.18 572.85 202.54 574.56 ;
   RECT 23.18 574.56 202.54 576.27 ;
   RECT 23.18 576.27 202.54 577.98 ;
   RECT 23.18 577.98 202.54 579.69 ;
   RECT 23.18 579.69 202.54 581.4 ;
   RECT 23.18 581.4 202.54 583.11 ;
   RECT 23.18 583.11 202.54 584.82 ;
   RECT 23.18 584.82 202.54 586.53 ;
   RECT 23.18 586.53 202.54 588.24 ;
   RECT 23.18 588.24 202.54 589.95 ;
   RECT 23.18 589.95 202.54 591.66 ;
   RECT 23.18 591.66 202.54 593.37 ;
   RECT 23.18 593.37 202.54 595.08 ;
   RECT 23.18 595.08 202.54 596.79 ;
   RECT 23.18 596.79 202.54 598.5 ;
   RECT 23.18 598.5 202.54 600.21 ;
   RECT 23.18 600.21 202.54 601.92 ;
   RECT 23.18 601.92 202.54 603.63 ;
   RECT 23.18 603.63 202.54 605.34 ;
   RECT 23.18 605.34 202.54 607.05 ;
   RECT 23.18 607.05 202.54 608.76 ;
   RECT 23.18 608.76 202.54 610.47 ;
   RECT 23.18 610.47 202.54 612.18 ;
   RECT 23.18 612.18 202.54 613.89 ;
   RECT 23.18 613.89 202.54 615.6 ;
   RECT 23.18 615.6 202.54 617.31 ;
   RECT 23.18 617.31 202.54 619.02 ;
   RECT 23.18 619.02 202.54 620.73 ;
   RECT 23.18 620.73 202.54 622.44 ;
   RECT 23.18 622.44 202.54 624.15 ;
   RECT 23.18 624.15 202.54 625.86 ;
   RECT 23.18 625.86 202.54 627.57 ;
   RECT 23.18 627.57 202.54 629.28 ;
   RECT 23.18 629.28 202.54 630.99 ;
   RECT 23.18 630.99 202.54 632.7 ;
   RECT 23.18 632.7 202.54 634.41 ;
   RECT 23.18 634.41 202.54 636.12 ;
   RECT 23.18 636.12 202.54 637.83 ;
   RECT 23.18 637.83 202.54 639.54 ;
   RECT 23.18 639.54 202.54 641.25 ;
   RECT 23.18 641.25 202.54 642.96 ;
   RECT 23.18 642.96 202.54 644.67 ;
   RECT 23.18 644.67 202.54 646.38 ;
   RECT 23.18 646.38 202.54 648.09 ;
   RECT 23.18 648.09 202.54 649.8 ;
   RECT 23.18 649.8 202.54 651.51 ;
   RECT 23.18 651.51 202.54 653.22 ;
   RECT 23.18 653.22 202.54 654.93 ;
   RECT 23.18 654.93 202.54 656.64 ;
   RECT 23.18 656.64 202.54 658.35 ;
   RECT 23.18 658.35 202.54 660.06 ;
   RECT 23.18 660.06 202.54 661.77 ;
   RECT 23.18 661.77 202.54 663.48 ;
   RECT 23.18 663.48 202.54 665.19 ;
   RECT 23.18 665.19 202.54 666.9 ;
   RECT 23.18 666.9 202.54 668.61 ;
   RECT 23.18 668.61 202.54 670.32 ;
   RECT 23.18 670.32 202.54 672.03 ;
   RECT 23.18 672.03 202.54 673.74 ;
   RECT 23.18 673.74 202.54 675.45 ;
   RECT 23.18 675.45 202.54 677.16 ;
   RECT 23.18 677.16 202.54 678.87 ;
   RECT 23.18 678.87 202.54 680.58 ;
   RECT 23.18 680.58 202.54 682.29 ;
   RECT 23.18 682.29 202.54 684.0 ;
   RECT 23.18 684.0 202.54 685.71 ;
   RECT 23.18 685.71 202.54 687.42 ;
   RECT 23.18 687.42 202.54 689.13 ;
   RECT 23.18 689.13 202.54 690.84 ;
   RECT 23.18 690.84 202.54 692.55 ;
   RECT 23.18 692.55 202.54 694.26 ;
   RECT 23.18 694.26 202.54 695.97 ;
   RECT 23.18 695.97 202.54 697.68 ;
   RECT 23.18 697.68 202.54 699.39 ;
   RECT 23.18 699.39 202.54 701.1 ;
   RECT 23.18 701.1 202.54 702.81 ;
   RECT 23.18 702.81 202.54 704.52 ;
   RECT 23.18 704.52 202.54 706.23 ;
   RECT 23.18 706.23 202.54 707.94 ;
   RECT 23.18 707.94 202.54 709.65 ;
   RECT 23.18 709.65 202.54 711.36 ;
   RECT 23.18 711.36 202.54 713.07 ;
   RECT 23.18 713.07 202.54 714.78 ;
   RECT 23.18 714.78 202.54 716.49 ;
   RECT 23.18 716.49 202.54 718.2 ;
   RECT 23.18 718.2 202.54 719.91 ;
   RECT 23.18 719.91 202.54 721.62 ;
   RECT 23.18 721.62 202.54 723.33 ;
   RECT 23.18 723.33 202.54 725.04 ;
   RECT 23.18 725.04 202.54 726.75 ;
   RECT 23.18 726.75 202.54 728.46 ;
   RECT 23.18 728.46 202.54 730.17 ;
   RECT 23.18 730.17 202.54 731.88 ;
   RECT 23.18 731.88 202.54 733.59 ;
   RECT 23.18 733.59 202.54 735.3 ;
   RECT 23.18 735.3 202.54 737.01 ;
   RECT 23.18 737.01 202.54 738.72 ;
   RECT 23.18 738.72 202.54 740.43 ;
   RECT 23.18 740.43 202.54 742.14 ;
   RECT 23.18 742.14 202.54 743.85 ;
   RECT 23.18 743.85 202.54 745.56 ;
   RECT 23.18 745.56 202.54 747.27 ;
   RECT 23.18 747.27 202.54 748.98 ;
   RECT 23.18 748.98 202.54 750.69 ;
   RECT 23.18 750.69 202.54 752.4 ;
   RECT 23.18 752.4 202.54 754.11 ;
   RECT 23.18 754.11 202.54 755.82 ;
   RECT 23.18 755.82 202.54 757.53 ;
   RECT 23.18 757.53 202.54 759.24 ;
   RECT 23.18 759.24 202.54 760.95 ;
   RECT 23.18 760.95 202.54 762.66 ;
   RECT 23.18 762.66 202.54 764.37 ;
   RECT 23.18 764.37 202.54 766.08 ;
   RECT 23.18 766.08 202.54 767.79 ;
   RECT 23.18 767.79 202.54 769.5 ;
   RECT 23.18 769.5 202.54 771.21 ;
   RECT 23.18 771.21 202.54 772.92 ;
   RECT 23.18 772.92 202.54 774.63 ;
   RECT 23.18 774.63 202.54 776.34 ;
   RECT 23.18 776.34 202.54 778.05 ;
   RECT 23.18 778.05 202.54 779.76 ;
   RECT 23.18 779.76 202.54 781.47 ;
   RECT 23.18 781.47 202.54 783.18 ;
   RECT 23.18 783.18 202.54 784.89 ;
   RECT 23.18 784.89 202.54 786.6 ;
   RECT 23.18 786.6 202.54 788.31 ;
   RECT 23.18 788.31 202.54 790.02 ;
   RECT 23.18 790.02 202.54 791.73 ;
   RECT 23.18 791.73 202.54 793.44 ;
   RECT 23.18 793.44 202.54 795.15 ;
   RECT 23.18 795.15 202.54 796.86 ;
   RECT 23.18 796.86 202.54 798.57 ;
   RECT 23.18 798.57 202.54 800.28 ;
   RECT 23.18 800.28 202.54 801.99 ;
   RECT 23.18 801.99 202.54 803.7 ;
   RECT 23.18 803.7 202.54 805.41 ;
   RECT 23.18 805.41 202.54 807.12 ;
   RECT 23.18 807.12 202.54 808.83 ;
   RECT 23.18 808.83 202.54 810.54 ;
   RECT 23.18 810.54 202.54 812.25 ;
   RECT 23.18 812.25 202.54 813.96 ;
   RECT 23.18 813.96 202.54 815.67 ;
   RECT 23.18 815.67 202.54 817.38 ;
   RECT 23.18 817.38 202.54 819.09 ;
   RECT 23.18 819.09 202.54 820.8 ;
   RECT 23.18 820.8 202.54 822.51 ;
   RECT 23.18 822.51 202.54 824.22 ;
   RECT 23.18 824.22 202.54 825.93 ;
   RECT 23.18 825.93 202.54 827.64 ;
   RECT 23.18 827.64 202.54 829.35 ;
   RECT 23.18 829.35 202.54 831.06 ;
   RECT 23.18 831.06 202.54 832.77 ;
   RECT 23.18 832.77 202.54 834.48 ;
   RECT 23.18 834.48 202.54 836.19 ;
   RECT 23.18 836.19 202.54 837.9 ;
   RECT 23.18 837.9 202.54 839.61 ;
   RECT 23.18 839.61 202.54 841.32 ;
 END
END block_533x4428_789

MACRO block_533x4428_789f
 CLASS BLOCK ;
 FOREIGN block_533x4428_789f 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 202.54 BY 841.32 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 834.96 176.22 835.52 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 830.77 176.22 831.35 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 794.11 176.22 794.67 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 360.71 176.22 361.29 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 356.54 176.22 357.11 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 352.55 176.22 353.12 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 348.37 176.22 348.94 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 344.38 176.22 344.94 ;
  END
 END o7
 PIN o8
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 340.19 176.22 340.76 ;
  END
 END o8
 PIN o9
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 336.20 176.22 336.77 ;
  END
 END o9
 PIN o10
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 332.02 176.22 332.60 ;
  END
 END o10
 PIN o11
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 328.04 176.22 328.61 ;
  END
 END o11
 PIN o12
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 323.86 176.22 324.43 ;
  END
 END o12
 PIN o13
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 789.92 176.22 790.50 ;
  END
 END o13
 PIN o14
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 319.87 176.22 320.44 ;
  END
 END o14
 PIN o15
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 315.69 176.22 316.25 ;
  END
 END o15
 PIN o16
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 293.45 176.22 294.02 ;
  END
 END o16
 PIN o17
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 289.27 176.22 289.85 ;
  END
 END o17
 PIN o18
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 285.29 176.22 285.86 ;
  END
 END o18
 PIN o19
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 281.11 176.22 281.68 ;
  END
 END o19
 PIN o20
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 277.12 176.22 277.69 ;
  END
 END o20
 PIN o21
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 272.94 176.22 273.50 ;
  END
 END o21
 PIN o22
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 268.94 176.22 269.51 ;
  END
 END o22
 PIN o23
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 264.76 176.22 265.33 ;
  END
 END o23
 PIN o24
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 785.93 176.22 786.50 ;
  END
 END o24
 PIN o25
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 260.77 176.22 261.35 ;
  END
 END o25
 PIN o26
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 256.60 176.22 257.17 ;
  END
 END o26
 PIN o27
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 252.60 176.22 253.18 ;
  END
 END o27
 PIN o28
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 248.43 176.22 249.00 ;
  END
 END o28
 PIN o29
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 244.44 176.22 245.00 ;
  END
 END o29
 PIN o30
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 240.25 176.22 240.82 ;
  END
 END o30
 PIN o31
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 236.26 176.22 236.84 ;
  END
 END o31
 PIN o32
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 232.09 176.22 232.66 ;
  END
 END o32
 PIN o33
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 228.09 176.22 228.66 ;
  END
 END o33
 PIN o34
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 223.91 176.22 224.49 ;
  END
 END o34
 PIN o35
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 781.75 176.22 782.33 ;
  END
 END o35
 PIN o36
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 219.93 176.22 220.50 ;
  END
 END o36
 PIN o37
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 215.75 176.22 216.31 ;
  END
 END o37
 PIN o38
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 211.75 176.22 212.32 ;
  END
 END o38
 PIN o39
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 207.57 176.22 208.15 ;
  END
 END o39
 PIN o40
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 198.46 176.22 199.03 ;
  END
 END o40
 PIN o41
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 194.28 176.22 194.84 ;
  END
 END o41
 PIN o42
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 190.28 176.22 190.85 ;
  END
 END o42
 PIN o43
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 186.10 176.22 186.68 ;
  END
 END o43
 PIN o44
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 182.12 176.22 182.69 ;
  END
 END o44
 PIN o45
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 177.94 176.22 178.50 ;
  END
 END o45
 PIN o46
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 777.76 176.22 778.34 ;
  END
 END o46
 PIN o47
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 173.94 176.22 174.51 ;
  END
 END o47
 PIN o48
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 169.76 176.22 170.34 ;
  END
 END o48
 PIN o49
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 165.78 176.22 166.34 ;
  END
 END o49
 PIN o50
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 161.59 176.22 162.16 ;
  END
 END o50
 PIN o51
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 157.60 176.22 158.18 ;
  END
 END o51
 PIN o52
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 153.43 176.22 154.00 ;
  END
 END o52
 PIN o53
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 149.44 176.22 150.00 ;
  END
 END o53
 PIN o54
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 145.25 176.22 145.82 ;
  END
 END o54
 PIN o55
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 141.26 176.22 141.84 ;
  END
 END o55
 PIN o56
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 137.09 176.22 137.66 ;
  END
 END o56
 PIN o57
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 773.59 176.22 774.15 ;
  END
 END o57
 PIN o58
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 133.09 176.22 133.66 ;
  END
 END o58
 PIN o59
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 128.91 176.22 129.49 ;
  END
 END o59
 PIN o60
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 124.92 176.22 125.50 ;
  END
 END o60
 PIN o61
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 120.75 176.22 121.31 ;
  END
 END o61
 PIN o62
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 116.75 176.22 117.33 ;
  END
 END o62
 PIN o63
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 112.58 176.22 113.14 ;
  END
 END o63
 PIN o64
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 90.34 176.22 90.92 ;
  END
 END o64
 PIN o65
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 86.17 176.22 86.73 ;
  END
 END o65
 PIN o66
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 82.17 176.22 82.75 ;
  END
 END o66
 PIN o67
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 78.00 176.22 78.56 ;
  END
 END o67
 PIN o68
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 769.60 176.22 770.16 ;
  END
 END o68
 PIN o69
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 74.00 176.22 74.58 ;
  END
 END o69
 PIN o70
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 69.83 176.22 70.39 ;
  END
 END o70
 PIN o71
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 65.83 176.22 66.41 ;
  END
 END o71
 PIN o72
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 61.66 176.22 62.23 ;
  END
 END o72
 PIN o73
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 57.66 176.22 58.23 ;
  END
 END o73
 PIN o74
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 53.48 176.22 54.05 ;
  END
 END o74
 PIN o75
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 49.49 176.22 50.06 ;
  END
 END o75
 PIN o76
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 45.31 176.22 45.88 ;
  END
 END o76
 PIN o77
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 41.33 176.22 41.90 ;
  END
 END o77
 PIN o78
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 37.15 176.22 37.72 ;
  END
 END o78
 PIN o79
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 765.41 176.22 765.99 ;
  END
 END o79
 PIN o80
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 33.16 176.22 33.73 ;
  END
 END o80
 PIN o81
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 28.98 176.22 29.55 ;
  END
 END o81
 PIN o82
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 24.98 176.22 25.55 ;
  END
 END o82
 PIN o83
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 20.80 176.22 21.38 ;
  END
 END o83
 PIN o84
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 16.82 176.22 17.39 ;
  END
 END o84
 PIN o85
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 12.63 176.22 13.21 ;
  END
 END o85
 PIN o86
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 8.64 176.22 9.21 ;
  END
 END o86
 PIN o87
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 4.46 176.22 5.04 ;
  END
 END o87
 PIN o88
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 761.42 176.22 762.00 ;
  END
 END o88
 PIN o89
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 757.25 176.22 757.82 ;
  END
 END o89
 PIN o90
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 826.78 176.22 827.36 ;
  END
 END o90
 PIN o91
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 753.25 176.22 753.83 ;
  END
 END o91
 PIN o92
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 749.08 176.22 749.64 ;
  END
 END o92
 PIN o93
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 745.09 176.22 745.65 ;
  END
 END o93
 PIN o94
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 722.66 176.22 723.24 ;
  END
 END o94
 PIN o95
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 718.67 176.22 719.25 ;
  END
 END o95
 PIN o96
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 714.50 176.22 715.07 ;
  END
 END o96
 PIN o97
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 710.50 176.22 711.08 ;
  END
 END o97
 PIN o98
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 706.33 176.22 706.89 ;
  END
 END o98
 PIN o99
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 702.34 176.22 702.90 ;
  END
 END o99
 PIN o100
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 698.15 176.22 698.73 ;
  END
 END o100
 PIN o101
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 822.61 176.22 823.17 ;
  END
 END o101
 PIN o102
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 694.16 176.22 694.74 ;
  END
 END o102
 PIN o103
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 689.99 176.22 690.55 ;
  END
 END o103
 PIN o104
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 686.00 176.22 686.57 ;
  END
 END o104
 PIN o105
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 681.82 176.22 682.38 ;
  END
 END o105
 PIN o106
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 677.83 176.22 678.39 ;
  END
 END o106
 PIN o107
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 673.64 176.22 674.22 ;
  END
 END o107
 PIN o108
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 669.65 176.22 670.23 ;
  END
 END o108
 PIN o109
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 665.48 176.22 666.04 ;
  END
 END o109
 PIN o110
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 661.49 176.22 662.05 ;
  END
 END o110
 PIN o111
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 657.30 176.22 657.88 ;
  END
 END o111
 PIN o112
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 818.62 176.22 819.18 ;
  END
 END o112
 PIN o113
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 653.32 176.22 653.88 ;
  END
 END o113
 PIN o114
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 649.13 176.22 649.71 ;
  END
 END o114
 PIN o115
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 645.14 176.22 645.72 ;
  END
 END o115
 PIN o116
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 640.97 176.22 641.53 ;
  END
 END o116
 PIN o117
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 636.98 176.22 637.54 ;
  END
 END o117
 PIN o118
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 632.79 176.22 633.37 ;
  END
 END o118
 PIN o119
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 623.67 176.22 624.25 ;
  END
 END o119
 PIN o120
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 619.50 176.22 620.07 ;
  END
 END o120
 PIN o121
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 615.50 176.22 616.08 ;
  END
 END o121
 PIN o122
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 611.33 176.22 611.89 ;
  END
 END o122
 PIN o123
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 814.43 176.22 815.00 ;
  END
 END o123
 PIN o124
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 607.34 176.22 607.90 ;
  END
 END o124
 PIN o125
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 603.15 176.22 603.73 ;
  END
 END o125
 PIN o126
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 599.16 176.22 599.74 ;
  END
 END o126
 PIN o127
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 594.99 176.22 595.55 ;
  END
 END o127
 PIN o128
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 591.00 176.22 591.57 ;
  END
 END o128
 PIN o129
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 586.82 176.22 587.38 ;
  END
 END o129
 PIN o130
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 582.83 176.22 583.39 ;
  END
 END o130
 PIN o131
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 578.64 176.22 579.22 ;
  END
 END o131
 PIN o132
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 574.65 176.22 575.23 ;
  END
 END o132
 PIN o133
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 570.48 176.22 571.04 ;
  END
 END o133
 PIN o134
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 810.45 176.22 811.01 ;
  END
 END o134
 PIN o135
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 566.49 176.22 567.05 ;
  END
 END o135
 PIN o136
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 562.30 176.22 562.88 ;
  END
 END o136
 PIN o137
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 558.32 176.22 558.88 ;
  END
 END o137
 PIN o138
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 554.13 176.22 554.71 ;
  END
 END o138
 PIN o139
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 550.14 176.22 550.72 ;
  END
 END o139
 PIN o140
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 545.97 176.22 546.53 ;
  END
 END o140
 PIN o141
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 541.98 176.22 542.54 ;
  END
 END o141
 PIN o142
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 537.79 176.22 538.37 ;
  END
 END o142
 PIN o143
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 515.57 176.22 516.13 ;
  END
 END o143
 PIN o144
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 511.38 176.22 511.95 ;
  END
 END o144
 PIN o145
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 806.26 176.22 806.84 ;
  END
 END o145
 PIN o146
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 507.39 176.22 507.96 ;
  END
 END o146
 PIN o147
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 503.21 176.22 503.79 ;
  END
 END o147
 PIN o148
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 499.23 176.22 499.80 ;
  END
 END o148
 PIN o149
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 495.05 176.22 495.62 ;
  END
 END o149
 PIN o150
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 491.06 176.22 491.62 ;
  END
 END o150
 PIN o151
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 486.88 176.22 487.44 ;
  END
 END o151
 PIN o152
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 482.88 176.22 483.45 ;
  END
 END o152
 PIN o153
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 478.70 176.22 479.27 ;
  END
 END o153
 PIN o154
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 474.71 176.22 475.29 ;
  END
 END o154
 PIN o155
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 470.54 176.22 471.11 ;
  END
 END o155
 PIN o156
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 802.27 176.22 802.85 ;
  END
 END o156
 PIN o157
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 466.55 176.22 467.12 ;
  END
 END o157
 PIN o158
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 462.37 176.22 462.94 ;
  END
 END o158
 PIN o159
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 458.38 176.22 458.94 ;
  END
 END o159
 PIN o160
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 454.19 176.22 454.76 ;
  END
 END o160
 PIN o161
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 450.20 176.22 450.77 ;
  END
 END o161
 PIN o162
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 446.02 176.22 446.60 ;
  END
 END o162
 PIN o163
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 442.04 176.22 442.61 ;
  END
 END o163
 PIN o164
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 437.86 176.22 438.43 ;
  END
 END o164
 PIN o165
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 433.87 176.22 434.44 ;
  END
 END o165
 PIN o166
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 429.69 176.22 430.25 ;
  END
 END o166
 PIN o167
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 798.10 176.22 798.66 ;
  END
 END o167
 PIN o168
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 401.56 176.22 402.13 ;
  END
 END o168
 PIN o169
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 397.38 176.22 397.95 ;
  END
 END o169
 PIN o170
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 393.39 176.22 393.96 ;
  END
 END o170
 PIN o171
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 389.21 176.22 389.79 ;
  END
 END o171
 PIN o172
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 385.23 176.22 385.80 ;
  END
 END o172
 PIN o173
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 381.05 176.22 381.62 ;
  END
 END o173
 PIN o174
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 377.06 176.22 377.62 ;
  END
 END o174
 PIN o175
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 372.88 176.22 373.44 ;
  END
 END o175
 PIN o176
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 368.88 176.22 369.45 ;
  END
 END o176
 PIN o177
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 364.70 176.22 365.27 ;
  END
 END o177
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.83 426.83 199.41 427.40 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.83 409.74 199.41 410.31 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.83 421.51 199.41 422.08 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.07 426.45 198.64 427.02 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.07 427.21 198.64 427.79 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.83 427.60 199.41 428.17 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.83 417.90 199.41 418.48 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.83 404.80 199.41 405.37 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.07 410.12 198.64 410.69 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.83 410.50 199.41 411.06 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.83 408.40 199.41 408.98 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.83 405.94 199.41 406.50 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.07 404.42 198.64 404.99 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 188.95 427.98 189.52 428.55 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 188.95 414.68 189.52 415.25 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 836.66 176.22 837.24 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 832.49 176.22 833.05 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 795.82 176.22 796.38 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 359.00 176.22 359.57 ;
  END
 END i18
 PIN i19
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 354.82 176.22 355.39 ;
  END
 END i19
 PIN i20
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 350.83 176.22 351.40 ;
  END
 END i20
 PIN i21
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 346.65 176.22 347.23 ;
  END
 END i21
 PIN i22
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 342.67 176.22 343.24 ;
  END
 END i22
 PIN i23
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 338.49 176.22 339.06 ;
  END
 END i23
 PIN i24
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 334.50 176.22 335.06 ;
  END
 END i24
 PIN i25
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 330.31 176.22 330.88 ;
  END
 END i25
 PIN i26
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 326.32 176.22 326.89 ;
  END
 END i26
 PIN i27
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 322.14 176.22 322.71 ;
  END
 END i27
 PIN i28
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 791.63 176.22 792.21 ;
  END
 END i28
 PIN i29
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 318.15 176.22 318.73 ;
  END
 END i29
 PIN i30
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 313.98 176.22 314.55 ;
  END
 END i30
 PIN i31
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 291.75 176.22 292.31 ;
  END
 END i31
 PIN i32
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 287.56 176.22 288.13 ;
  END
 END i32
 PIN i33
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 283.57 176.22 284.14 ;
  END
 END i33
 PIN i34
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 279.39 176.22 279.96 ;
  END
 END i34
 PIN i35
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 275.40 176.22 275.98 ;
  END
 END i35
 PIN i36
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 271.23 176.22 271.80 ;
  END
 END i36
 PIN i37
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 267.24 176.22 267.81 ;
  END
 END i37
 PIN i38
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 263.06 176.22 263.62 ;
  END
 END i38
 PIN i39
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 787.64 176.22 788.22 ;
  END
 END i39
 PIN i40
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 259.06 176.22 259.63 ;
  END
 END i40
 PIN i41
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 254.88 176.22 255.46 ;
  END
 END i41
 PIN i42
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 250.90 176.22 251.47 ;
  END
 END i42
 PIN i43
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 246.72 176.22 247.28 ;
  END
 END i43
 PIN i44
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 242.72 176.22 243.29 ;
  END
 END i44
 PIN i45
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 238.54 176.22 239.12 ;
  END
 END i45
 PIN i46
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 234.56 176.22 235.12 ;
  END
 END i46
 PIN i47
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 230.38 176.22 230.94 ;
  END
 END i47
 PIN i48
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 226.38 176.22 226.96 ;
  END
 END i48
 PIN i49
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 222.21 176.22 222.78 ;
  END
 END i49
 PIN i50
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 783.47 176.22 784.03 ;
  END
 END i50
 PIN i51
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 218.22 176.22 218.78 ;
  END
 END i51
 PIN i52
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 214.03 176.22 214.60 ;
  END
 END i52
 PIN i53
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 210.04 176.22 210.62 ;
  END
 END i53
 PIN i54
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 205.87 176.22 206.44 ;
  END
 END i54
 PIN i55
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 196.75 176.22 197.31 ;
  END
 END i55
 PIN i56
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 192.56 176.22 193.13 ;
  END
 END i56
 PIN i57
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 188.57 176.22 189.15 ;
  END
 END i57
 PIN i58
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 184.40 176.22 184.97 ;
  END
 END i58
 PIN i59
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 180.41 176.22 180.97 ;
  END
 END i59
 PIN i60
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 176.22 176.22 176.79 ;
  END
 END i60
 PIN i61
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 779.48 176.22 780.04 ;
  END
 END i61
 PIN i62
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 172.24 176.22 172.81 ;
  END
 END i62
 PIN i63
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 168.06 176.22 168.62 ;
  END
 END i63
 PIN i64
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 164.06 176.22 164.63 ;
  END
 END i64
 PIN i65
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 159.88 176.22 160.46 ;
  END
 END i65
 PIN i66
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 155.90 176.22 156.47 ;
  END
 END i66
 PIN i67
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 151.72 176.22 152.28 ;
  END
 END i67
 PIN i68
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 147.72 176.22 148.29 ;
  END
 END i68
 PIN i69
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 143.54 176.22 144.12 ;
  END
 END i69
 PIN i70
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 139.56 176.22 140.12 ;
  END
 END i70
 PIN i71
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 135.38 176.22 135.94 ;
  END
 END i71
 PIN i72
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 775.29 176.22 775.87 ;
  END
 END i72
 PIN i73
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 131.38 176.22 131.96 ;
  END
 END i73
 PIN i74
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 127.20 176.22 127.78 ;
  END
 END i74
 PIN i75
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 123.22 176.22 123.78 ;
  END
 END i75
 PIN i76
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 119.03 176.22 119.61 ;
  END
 END i76
 PIN i77
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 115.05 176.22 115.61 ;
  END
 END i77
 PIN i78
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 110.86 176.22 111.44 ;
  END
 END i78
 PIN i79
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 88.64 176.22 89.20 ;
  END
 END i79
 PIN i80
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 84.45 176.22 85.03 ;
  END
 END i80
 PIN i81
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 80.47 176.22 81.03 ;
  END
 END i81
 PIN i82
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 76.28 176.22 76.86 ;
  END
 END i82
 PIN i83
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 771.30 176.22 771.88 ;
  END
 END i83
 PIN i84
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 72.30 176.22 72.86 ;
  END
 END i84
 PIN i85
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 68.11 176.22 68.69 ;
  END
 END i85
 PIN i86
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 64.12 176.22 64.69 ;
  END
 END i86
 PIN i87
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 59.95 176.22 60.52 ;
  END
 END i87
 PIN i88
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 55.95 176.22 56.52 ;
  END
 END i88
 PIN i89
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 51.77 176.22 52.34 ;
  END
 END i89
 PIN i90
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 47.78 176.22 48.35 ;
  END
 END i90
 PIN i91
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 43.60 176.22 44.17 ;
  END
 END i91
 PIN i92
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 39.62 176.22 40.19 ;
  END
 END i92
 PIN i93
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 35.44 176.22 36.01 ;
  END
 END i93
 PIN i94
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 767.12 176.22 767.70 ;
  END
 END i94
 PIN i95
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 31.45 176.22 32.02 ;
  END
 END i95
 PIN i96
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 27.27 176.22 27.84 ;
  END
 END i96
 PIN i97
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 23.27 176.22 23.84 ;
  END
 END i97
 PIN i98
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 19.09 176.22 19.66 ;
  END
 END i98
 PIN i99
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 15.11 176.22 15.68 ;
  END
 END i99
 PIN i100
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 10.93 176.22 11.49 ;
  END
 END i100
 PIN i101
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 6.93 176.22 7.50 ;
  END
 END i101
 PIN i102
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 2.75 176.22 3.33 ;
  END
 END i102
 PIN i103
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 763.13 176.22 763.71 ;
  END
 END i103
 PIN i104
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 758.96 176.22 759.52 ;
  END
 END i104
 PIN i105
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 828.50 176.22 829.07 ;
  END
 END i105
 PIN i106
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 754.97 176.22 755.53 ;
  END
 END i106
 PIN i107
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 750.78 176.22 751.36 ;
  END
 END i107
 PIN i108
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 746.79 176.22 747.37 ;
  END
 END i108
 PIN i109
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 724.38 176.22 724.95 ;
  END
 END i109
 PIN i110
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 720.38 176.22 720.96 ;
  END
 END i110
 PIN i111
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 716.21 176.22 716.77 ;
  END
 END i111
 PIN i112
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 712.22 176.22 712.78 ;
  END
 END i112
 PIN i113
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 708.03 176.22 708.61 ;
  END
 END i113
 PIN i114
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 704.04 176.22 704.62 ;
  END
 END i114
 PIN i115
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 699.87 176.22 700.43 ;
  END
 END i115
 PIN i116
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 824.32 176.22 824.88 ;
  END
 END i116
 PIN i117
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 695.88 176.22 696.45 ;
  END
 END i117
 PIN i118
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 691.70 176.22 692.26 ;
  END
 END i118
 PIN i119
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 687.71 176.22 688.27 ;
  END
 END i119
 PIN i120
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 683.52 176.22 684.10 ;
  END
 END i120
 PIN i121
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 679.53 176.22 680.11 ;
  END
 END i121
 PIN i122
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 675.36 176.22 675.92 ;
  END
 END i122
 PIN i123
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 671.37 176.22 671.93 ;
  END
 END i123
 PIN i124
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 667.18 176.22 667.75 ;
  END
 END i124
 PIN i125
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 663.20 176.22 663.76 ;
  END
 END i125
 PIN i126
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 659.01 176.22 659.59 ;
  END
 END i126
 PIN i127
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 820.33 176.22 820.89 ;
  END
 END i127
 PIN i128
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 655.02 176.22 655.60 ;
  END
 END i128
 PIN i129
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 650.85 176.22 651.41 ;
  END
 END i129
 PIN i130
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 646.86 176.22 647.42 ;
  END
 END i130
 PIN i131
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 642.67 176.22 643.25 ;
  END
 END i131
 PIN i132
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 638.68 176.22 639.25 ;
  END
 END i132
 PIN i133
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 634.50 176.22 635.08 ;
  END
 END i133
 PIN i134
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 625.38 176.22 625.96 ;
  END
 END i134
 PIN i135
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 621.21 176.22 621.77 ;
  END
 END i135
 PIN i136
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 617.22 176.22 617.78 ;
  END
 END i136
 PIN i137
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 613.03 176.22 613.61 ;
  END
 END i137
 PIN i138
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 816.14 176.22 816.72 ;
  END
 END i138
 PIN i139
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 609.04 176.22 609.62 ;
  END
 END i139
 PIN i140
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 604.87 176.22 605.43 ;
  END
 END i140
 PIN i141
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 600.88 176.22 601.45 ;
  END
 END i141
 PIN i142
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 596.70 176.22 597.26 ;
  END
 END i142
 PIN i143
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 592.71 176.22 593.27 ;
  END
 END i143
 PIN i144
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 588.52 176.22 589.10 ;
  END
 END i144
 PIN i145
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 584.53 176.22 585.11 ;
  END
 END i145
 PIN i146
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 580.36 176.22 580.92 ;
  END
 END i146
 PIN i147
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 576.37 176.22 576.93 ;
  END
 END i147
 PIN i148
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 572.18 176.22 572.75 ;
  END
 END i148
 PIN i149
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 812.15 176.22 812.73 ;
  END
 END i149
 PIN i150
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 568.20 176.22 568.76 ;
  END
 END i150
 PIN i151
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 564.01 176.22 564.59 ;
  END
 END i151
 PIN i152
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 560.02 176.22 560.60 ;
  END
 END i152
 PIN i153
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 555.85 176.22 556.41 ;
  END
 END i153
 PIN i154
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 551.86 176.22 552.42 ;
  END
 END i154
 PIN i155
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 547.67 176.22 548.25 ;
  END
 END i155
 PIN i156
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 543.68 176.22 544.25 ;
  END
 END i156
 PIN i157
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 539.50 176.22 540.08 ;
  END
 END i157
 PIN i158
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 517.27 176.22 517.85 ;
  END
 END i158
 PIN i159
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 513.10 176.22 513.66 ;
  END
 END i159
 PIN i160
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 807.98 176.22 808.54 ;
  END
 END i160
 PIN i161
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 509.11 176.22 509.68 ;
  END
 END i161
 PIN i162
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 504.93 176.22 505.50 ;
  END
 END i162
 PIN i163
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 500.94 176.22 501.50 ;
  END
 END i163
 PIN i164
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 496.75 176.22 497.32 ;
  END
 END i164
 PIN i165
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 492.76 176.22 493.33 ;
  END
 END i165
 PIN i166
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 488.58 176.22 489.15 ;
  END
 END i166
 PIN i167
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 484.60 176.22 485.17 ;
  END
 END i167
 PIN i168
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 480.42 176.22 480.99 ;
  END
 END i168
 PIN i169
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 476.43 176.22 477.00 ;
  END
 END i169
 PIN i170
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 472.25 176.22 472.81 ;
  END
 END i170
 PIN i171
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 803.99 176.22 804.55 ;
  END
 END i171
 PIN i172
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 468.25 176.22 468.82 ;
  END
 END i172
 PIN i173
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 464.07 176.22 464.64 ;
  END
 END i173
 PIN i174
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 460.08 176.22 460.65 ;
  END
 END i174
 PIN i175
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 455.90 176.22 456.48 ;
  END
 END i175
 PIN i176
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 451.92 176.22 452.49 ;
  END
 END i176
 PIN i177
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 447.74 176.22 448.31 ;
  END
 END i177
 PIN i178
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 443.75 176.22 444.31 ;
  END
 END i178
 PIN i179
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 439.56 176.22 440.13 ;
  END
 END i179
 PIN i180
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 435.57 176.22 436.14 ;
  END
 END i180
 PIN i181
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 431.39 176.22 431.96 ;
  END
 END i181
 PIN i182
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 799.80 176.22 800.38 ;
  END
 END i182
 PIN i183
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 399.86 176.22 400.43 ;
  END
 END i183
 PIN i184
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 395.68 176.22 396.25 ;
  END
 END i184
 PIN i185
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 391.69 176.22 392.25 ;
  END
 END i185
 PIN i186
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 387.50 176.22 388.07 ;
  END
 END i186
 PIN i187
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 383.51 176.22 384.08 ;
  END
 END i187
 PIN i188
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 379.33 176.22 379.90 ;
  END
 END i188
 PIN i189
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 375.35 176.22 375.92 ;
  END
 END i189
 PIN i190
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 371.17 176.22 371.74 ;
  END
 END i190
 PIN i191
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 367.18 176.22 367.75 ;
  END
 END i191
 PIN i192
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 175.66 363.00 176.22 363.56 ;
  END
 END i192
 PIN i193
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 769.02 175.47 769.60 ;
  END
 END i193
 PIN i194
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 764.85 175.47 765.41 ;
  END
 END i194
 PIN i195
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 760.86 175.47 761.42 ;
  END
 END i195
 PIN i196
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 781.18 175.47 781.75 ;
  END
 END i196
 PIN i197
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 777.20 175.47 777.76 ;
  END
 END i197
 PIN i198
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 701.76 175.47 702.34 ;
  END
 END i198
 PIN i199
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 697.59 175.47 698.15 ;
  END
 END i199
 PIN i200
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 693.60 175.47 694.16 ;
  END
 END i200
 PIN i201
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 689.41 175.47 689.99 ;
  END
 END i201
 PIN i202
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 685.42 175.47 686.00 ;
  END
 END i202
 PIN i203
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 561.74 175.47 562.30 ;
  END
 END i203
 PIN i204
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 557.75 175.47 558.32 ;
  END
 END i204
 PIN i205
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 553.57 175.47 554.13 ;
  END
 END i205
 PIN i206
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 574.09 175.47 574.65 ;
  END
 END i206
 PIN i207
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 569.90 175.47 570.48 ;
  END
 END i207
 PIN i208
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 494.48 175.47 495.05 ;
  END
 END i208
 PIN i209
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 490.49 175.47 491.06 ;
  END
 END i209
 PIN i210
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 486.31 175.47 486.88 ;
  END
 END i210
 PIN i211
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 482.31 175.47 482.88 ;
  END
 END i211
 PIN i212
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 478.13 175.47 478.70 ;
  END
 END i212
 PIN i213
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 336.77 175.47 337.35 ;
  END
 END i213
 PIN i214
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 340.76 175.47 341.33 ;
  END
 END i214
 PIN i215
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 344.94 175.47 345.51 ;
  END
 END i215
 PIN i216
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 348.94 175.47 349.50 ;
  END
 END i216
 PIN i217
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 353.12 175.47 353.69 ;
  END
 END i217
 PIN i218
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 269.51 175.47 270.08 ;
  END
 END i218
 PIN i219
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 273.50 175.47 274.07 ;
  END
 END i219
 PIN i220
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 277.69 175.47 278.25 ;
  END
 END i220
 PIN i221
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 257.17 175.47 257.74 ;
  END
 END i221
 PIN i222
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 261.35 175.47 261.92 ;
  END
 END i222
 PIN i223
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 133.66 175.47 134.24 ;
  END
 END i223
 PIN i224
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 137.66 175.47 138.22 ;
  END
 END i224
 PIN i225
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 141.84 175.47 142.41 ;
  END
 END i225
 PIN i226
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 145.82 175.47 146.40 ;
  END
 END i226
 PIN i227
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 150.00 175.47 150.57 ;
  END
 END i227
 PIN i228
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 66.41 175.47 66.97 ;
  END
 END i228
 PIN i229
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 70.39 175.47 70.97 ;
  END
 END i229
 PIN i230
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 74.58 175.47 75.14 ;
  END
 END i230
 PIN i231
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 54.05 175.47 54.62 ;
  END
 END i231
 PIN i232
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 58.23 175.47 58.80 ;
  END
 END i232
 PIN i233
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 773.01 175.47 773.59 ;
  END
 END i233
 PIN i234
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 705.75 175.47 706.33 ;
  END
 END i234
 PIN i235
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 565.91 175.47 566.49 ;
  END
 END i235
 PIN i236
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 498.65 175.47 499.23 ;
  END
 END i236
 PIN i237
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 332.60 175.47 333.17 ;
  END
 END i237
 PIN i238
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 265.33 175.47 265.90 ;
  END
 END i238
 PIN i239
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 129.49 175.47 130.06 ;
  END
 END i239
 PIN i240
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 62.23 175.47 62.80 ;
  END
 END i240
 PIN i241
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 184.01 427.98 184.58 428.55 ;
  END
 END i241
 PIN i242
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 184.01 414.68 184.58 415.25 ;
  END
 END i242
 PIN i243
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 836.10 175.47 836.66 ;
  END
 END i243
 PIN i244
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 831.91 175.47 832.49 ;
  END
 END i244
 PIN i245
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 795.25 175.47 795.82 ;
  END
 END i245
 PIN i246
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 359.57 175.47 360.14 ;
  END
 END i246
 PIN i247
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 355.39 175.47 355.96 ;
  END
 END i247
 PIN i248
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 351.40 175.47 351.98 ;
  END
 END i248
 PIN i249
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 347.23 175.47 347.80 ;
  END
 END i249
 PIN i250
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 343.24 175.47 343.81 ;
  END
 END i250
 PIN i251
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 339.06 175.47 339.62 ;
  END
 END i251
 PIN i252
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 335.06 175.47 335.63 ;
  END
 END i252
 PIN i253
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 330.88 175.47 331.45 ;
  END
 END i253
 PIN i254
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 326.89 175.47 327.46 ;
  END
 END i254
 PIN i255
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 322.71 175.47 323.29 ;
  END
 END i255
 PIN i256
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 791.07 175.47 791.63 ;
  END
 END i256
 PIN i257
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 318.73 175.47 319.30 ;
  END
 END i257
 PIN i258
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 314.55 175.47 315.12 ;
  END
 END i258
 PIN i259
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 292.31 175.47 292.88 ;
  END
 END i259
 PIN i260
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 288.13 175.47 288.70 ;
  END
 END i260
 PIN i261
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 284.14 175.47 284.71 ;
  END
 END i261
 PIN i262
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 279.96 175.47 280.54 ;
  END
 END i262
 PIN i263
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 275.98 175.47 276.55 ;
  END
 END i263
 PIN i264
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 271.80 175.47 272.37 ;
  END
 END i264
 PIN i265
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 267.81 175.47 268.38 ;
  END
 END i265
 PIN i266
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 263.62 175.47 264.19 ;
  END
 END i266
 PIN i267
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 787.08 175.47 787.64 ;
  END
 END i267
 PIN i268
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 259.63 175.47 260.20 ;
  END
 END i268
 PIN i269
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 255.46 175.47 256.02 ;
  END
 END i269
 PIN i270
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 251.47 175.47 252.03 ;
  END
 END i270
 PIN i271
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 247.28 175.47 247.85 ;
  END
 END i271
 PIN i272
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 243.29 175.47 243.87 ;
  END
 END i272
 PIN i273
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 239.12 175.47 239.69 ;
  END
 END i273
 PIN i274
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 235.12 175.47 235.69 ;
  END
 END i274
 PIN i275
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 230.94 175.47 231.51 ;
  END
 END i275
 PIN i276
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 226.96 175.47 227.53 ;
  END
 END i276
 PIN i277
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 222.78 175.47 223.34 ;
  END
 END i277
 PIN i278
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 782.89 175.47 783.47 ;
  END
 END i278
 PIN i279
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 218.78 175.47 219.35 ;
  END
 END i279
 PIN i280
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 214.60 175.47 215.18 ;
  END
 END i280
 PIN i281
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 210.62 175.47 211.19 ;
  END
 END i281
 PIN i282
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 206.44 175.47 207.00 ;
  END
 END i282
 PIN i283
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 197.31 175.47 197.88 ;
  END
 END i283
 PIN i284
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 193.13 175.47 193.71 ;
  END
 END i284
 PIN i285
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 189.15 175.47 189.72 ;
  END
 END i285
 PIN i286
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 184.97 175.47 185.53 ;
  END
 END i286
 PIN i287
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 180.97 175.47 181.54 ;
  END
 END i287
 PIN i288
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 176.79 175.47 177.37 ;
  END
 END i288
 PIN i289
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 778.90 175.47 779.48 ;
  END
 END i289
 PIN i290
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 172.81 175.47 173.38 ;
  END
 END i290
 PIN i291
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 168.62 175.47 169.19 ;
  END
 END i291
 PIN i292
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 164.63 175.47 165.21 ;
  END
 END i292
 PIN i293
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 160.46 175.47 161.03 ;
  END
 END i293
 PIN i294
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 156.47 175.47 157.03 ;
  END
 END i294
 PIN i295
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 152.28 175.47 152.85 ;
  END
 END i295
 PIN i296
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 148.29 175.47 148.87 ;
  END
 END i296
 PIN i297
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 144.12 175.47 144.69 ;
  END
 END i297
 PIN i298
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 140.12 175.47 140.69 ;
  END
 END i298
 PIN i299
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 135.94 175.47 136.51 ;
  END
 END i299
 PIN i300
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 774.73 175.47 775.29 ;
  END
 END i300
 PIN i301
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 131.96 175.47 132.53 ;
  END
 END i301
 PIN i302
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 127.78 175.47 128.34 ;
  END
 END i302
 PIN i303
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 123.78 175.47 124.36 ;
  END
 END i303
 PIN i304
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 119.61 175.47 120.17 ;
  END
 END i304
 PIN i305
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 115.61 175.47 116.19 ;
  END
 END i305
 PIN i306
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 111.44 175.47 112.00 ;
  END
 END i306
 PIN i307
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 89.20 175.47 89.78 ;
  END
 END i307
 PIN i308
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 85.03 175.47 85.59 ;
  END
 END i308
 PIN i309
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 81.03 175.47 81.61 ;
  END
 END i309
 PIN i310
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 76.86 175.47 77.42 ;
  END
 END i310
 PIN i311
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 770.74 175.47 771.30 ;
  END
 END i311
 PIN i312
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 72.86 175.47 73.44 ;
  END
 END i312
 PIN i313
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 68.69 175.47 69.25 ;
  END
 END i313
 PIN i314
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 64.69 175.47 65.27 ;
  END
 END i314
 PIN i315
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 60.52 175.47 61.09 ;
  END
 END i315
 PIN i316
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 56.52 175.47 57.09 ;
  END
 END i316
 PIN i317
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 52.34 175.47 52.91 ;
  END
 END i317
 PIN i318
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 48.35 175.47 48.92 ;
  END
 END i318
 PIN i319
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 44.17 175.47 44.74 ;
  END
 END i319
 PIN i320
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 40.19 175.47 40.76 ;
  END
 END i320
 PIN i321
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 36.01 175.47 36.58 ;
  END
 END i321
 PIN i322
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 766.55 175.47 767.12 ;
  END
 END i322
 PIN i323
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 32.02 175.47 32.59 ;
  END
 END i323
 PIN i324
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 27.84 175.47 28.41 ;
  END
 END i324
 PIN i325
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 23.84 175.47 24.41 ;
  END
 END i325
 PIN i326
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 19.66 175.47 20.23 ;
  END
 END i326
 PIN i327
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 15.68 175.47 16.25 ;
  END
 END i327
 PIN i328
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 11.49 175.47 12.06 ;
  END
 END i328
 PIN i329
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 7.50 175.47 8.07 ;
  END
 END i329
 PIN i330
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 3.33 175.47 3.90 ;
  END
 END i330
 PIN i331
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 762.57 175.47 763.13 ;
  END
 END i331
 PIN i332
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 758.38 175.47 758.96 ;
  END
 END i332
 PIN i333
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 827.92 175.47 828.50 ;
  END
 END i333
 PIN i334
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 754.39 175.47 754.97 ;
  END
 END i334
 PIN i335
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 750.22 175.47 750.78 ;
  END
 END i335
 PIN i336
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 746.23 175.47 746.79 ;
  END
 END i336
 PIN i337
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 723.80 175.47 724.38 ;
  END
 END i337
 PIN i338
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 719.82 175.47 720.38 ;
  END
 END i338
 PIN i339
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 715.63 175.47 716.21 ;
  END
 END i339
 PIN i340
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 711.64 175.47 712.22 ;
  END
 END i340
 PIN i341
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 707.47 175.47 708.03 ;
  END
 END i341
 PIN i342
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 703.48 175.47 704.04 ;
  END
 END i342
 PIN i343
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 699.29 175.47 699.87 ;
  END
 END i343
 PIN i344
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 823.75 175.47 824.32 ;
  END
 END i344
 PIN i345
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 695.30 175.47 695.88 ;
  END
 END i345
 PIN i346
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 691.12 175.47 691.70 ;
  END
 END i346
 PIN i347
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 687.13 175.47 687.71 ;
  END
 END i347
 PIN i348
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 682.96 175.47 683.52 ;
  END
 END i348
 PIN i349
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 678.97 175.47 679.53 ;
  END
 END i349
 PIN i350
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 674.78 175.47 675.36 ;
  END
 END i350
 PIN i351
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 670.79 175.47 671.37 ;
  END
 END i351
 PIN i352
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 666.62 175.47 667.18 ;
  END
 END i352
 PIN i353
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 662.62 175.47 663.20 ;
  END
 END i353
 PIN i354
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 658.45 175.47 659.01 ;
  END
 END i354
 PIN i355
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 819.75 175.47 820.33 ;
  END
 END i355
 PIN i356
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 654.46 175.47 655.02 ;
  END
 END i356
 PIN i357
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 650.27 175.47 650.85 ;
  END
 END i357
 PIN i358
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 646.28 175.47 646.86 ;
  END
 END i358
 PIN i359
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 642.11 175.47 642.67 ;
  END
 END i359
 PIN i360
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 638.12 175.47 638.68 ;
  END
 END i360
 PIN i361
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 633.93 175.47 634.50 ;
  END
 END i361
 PIN i362
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 624.82 175.47 625.38 ;
  END
 END i362
 PIN i363
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 620.63 175.47 621.21 ;
  END
 END i363
 PIN i364
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 616.64 175.47 617.22 ;
  END
 END i364
 PIN i365
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 612.47 175.47 613.03 ;
  END
 END i365
 PIN i366
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 815.58 175.47 816.14 ;
  END
 END i366
 PIN i367
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 608.48 175.47 609.04 ;
  END
 END i367
 PIN i368
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 604.29 175.47 604.87 ;
  END
 END i368
 PIN i369
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 600.30 175.47 600.88 ;
  END
 END i369
 PIN i370
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 596.12 175.47 596.70 ;
  END
 END i370
 PIN i371
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 592.13 175.47 592.71 ;
  END
 END i371
 PIN i372
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 587.96 175.47 588.52 ;
  END
 END i372
 PIN i373
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 583.97 175.47 584.53 ;
  END
 END i373
 PIN i374
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 579.78 175.47 580.36 ;
  END
 END i374
 PIN i375
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 575.79 175.47 576.37 ;
  END
 END i375
 PIN i376
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 571.62 175.47 572.18 ;
  END
 END i376
 PIN i377
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 811.59 175.47 812.15 ;
  END
 END i377
 PIN i378
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 567.62 175.47 568.20 ;
  END
 END i378
 PIN i379
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 563.45 175.47 564.01 ;
  END
 END i379
 PIN i380
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 559.46 175.47 560.02 ;
  END
 END i380
 PIN i381
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 555.27 175.47 555.85 ;
  END
 END i381
 PIN i382
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 551.28 175.47 551.86 ;
  END
 END i382
 PIN i383
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 547.11 175.47 547.67 ;
  END
 END i383
 PIN i384
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 543.12 175.47 543.68 ;
  END
 END i384
 PIN i385
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 538.93 175.47 539.50 ;
  END
 END i385
 PIN i386
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 516.71 175.47 517.27 ;
  END
 END i386
 PIN i387
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 512.52 175.47 513.10 ;
  END
 END i387
 PIN i388
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 807.40 175.47 807.98 ;
  END
 END i388
 PIN i389
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 508.54 175.47 509.11 ;
  END
 END i389
 PIN i390
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 504.36 175.47 504.93 ;
  END
 END i390
 PIN i391
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 500.37 175.47 500.94 ;
  END
 END i391
 PIN i392
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 496.19 175.47 496.75 ;
  END
 END i392
 PIN i393
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 492.19 175.47 492.76 ;
  END
 END i393
 PIN i394
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 488.01 175.47 488.58 ;
  END
 END i394
 PIN i395
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 484.02 175.47 484.60 ;
  END
 END i395
 PIN i396
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 479.85 175.47 480.42 ;
  END
 END i396
 PIN i397
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 475.86 175.47 476.43 ;
  END
 END i397
 PIN i398
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 471.68 175.47 472.25 ;
  END
 END i398
 PIN i399
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 803.41 175.47 803.99 ;
  END
 END i399
 PIN i400
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 467.69 175.47 468.25 ;
  END
 END i400
 PIN i401
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 463.50 175.47 464.07 ;
  END
 END i401
 PIN i402
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 459.51 175.47 460.08 ;
  END
 END i402
 PIN i403
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 455.33 175.47 455.90 ;
  END
 END i403
 PIN i404
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 451.35 175.47 451.92 ;
  END
 END i404
 PIN i405
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 447.17 175.47 447.74 ;
  END
 END i405
 PIN i406
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 443.18 175.47 443.75 ;
  END
 END i406
 PIN i407
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 439.00 175.47 439.56 ;
  END
 END i407
 PIN i408
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 435.00 175.47 435.57 ;
  END
 END i408
 PIN i409
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 430.82 175.47 431.39 ;
  END
 END i409
 PIN i410
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 799.24 175.47 799.80 ;
  END
 END i410
 PIN i411
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 400.43 175.47 401.00 ;
  END
 END i411
 PIN i412
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 396.25 175.47 396.81 ;
  END
 END i412
 PIN i413
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 392.25 175.47 392.82 ;
  END
 END i413
 PIN i414
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 388.07 175.47 388.64 ;
  END
 END i414
 PIN i415
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 384.08 175.47 384.65 ;
  END
 END i415
 PIN i416
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 379.90 175.47 380.48 ;
  END
 END i416
 PIN i417
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 375.92 175.47 376.49 ;
  END
 END i417
 PIN i418
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 371.74 175.47 372.31 ;
  END
 END i418
 PIN i419
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 367.75 175.47 368.31 ;
  END
 END i419
 PIN i420
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.89 363.56 175.47 364.13 ;
  END
 END i420
 PIN i421
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.83 420.38 199.41 420.94 ;
  END
 END i421
 PIN i422
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 198.07 420.00 198.64 420.56 ;
  END
 END i422
 PIN i423
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 835.52 174.70 836.10 ;
  END
 END i423
 PIN i424
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 831.35 174.70 831.91 ;
  END
 END i424
 PIN i425
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 794.67 174.70 795.25 ;
  END
 END i425
 PIN i426
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 360.14 174.70 360.71 ;
  END
 END i426
 PIN i427
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 355.96 174.70 356.54 ;
  END
 END i427
 PIN i428
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 351.98 174.70 352.55 ;
  END
 END i428
 PIN i429
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 347.80 174.70 348.37 ;
  END
 END i429
 PIN i430
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 343.81 174.70 344.38 ;
  END
 END i430
 PIN i431
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 339.62 174.70 340.19 ;
  END
 END i431
 PIN i432
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 335.63 174.70 336.20 ;
  END
 END i432
 PIN i433
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 331.45 174.70 332.02 ;
  END
 END i433
 PIN i434
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 327.46 174.70 328.04 ;
  END
 END i434
 PIN i435
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 323.29 174.70 323.86 ;
  END
 END i435
 PIN i436
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 790.50 174.70 791.07 ;
  END
 END i436
 PIN i437
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 319.30 174.70 319.87 ;
  END
 END i437
 PIN i438
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 315.12 174.70 315.69 ;
  END
 END i438
 PIN i439
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 292.88 174.70 293.45 ;
  END
 END i439
 PIN i440
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 288.70 174.70 289.27 ;
  END
 END i440
 PIN i441
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 284.71 174.70 285.29 ;
  END
 END i441
 PIN i442
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 280.54 174.70 281.11 ;
  END
 END i442
 PIN i443
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 276.55 174.70 277.12 ;
  END
 END i443
 PIN i444
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 272.37 174.70 272.94 ;
  END
 END i444
 PIN i445
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 268.38 174.70 268.94 ;
  END
 END i445
 PIN i446
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 264.19 174.70 264.76 ;
  END
 END i446
 PIN i447
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 786.50 174.70 787.08 ;
  END
 END i447
 PIN i448
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 260.20 174.70 260.77 ;
  END
 END i448
 PIN i449
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 256.02 174.70 256.60 ;
  END
 END i449
 PIN i450
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 252.03 174.70 252.60 ;
  END
 END i450
 PIN i451
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 247.85 174.70 248.43 ;
  END
 END i451
 PIN i452
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 243.87 174.70 244.44 ;
  END
 END i452
 PIN i453
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 239.69 174.70 240.25 ;
  END
 END i453
 PIN i454
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 235.69 174.70 236.26 ;
  END
 END i454
 PIN i455
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 231.51 174.70 232.09 ;
  END
 END i455
 PIN i456
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 227.53 174.70 228.09 ;
  END
 END i456
 PIN i457
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 223.34 174.70 223.91 ;
  END
 END i457
 PIN i458
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 782.33 174.70 782.89 ;
  END
 END i458
 PIN i459
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 219.35 174.70 219.93 ;
  END
 END i459
 PIN i460
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 215.18 174.70 215.75 ;
  END
 END i460
 PIN i461
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 211.19 174.70 211.75 ;
  END
 END i461
 PIN i462
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 207.00 174.70 207.57 ;
  END
 END i462
 PIN i463
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 197.88 174.70 198.46 ;
  END
 END i463
 PIN i464
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 193.71 174.70 194.28 ;
  END
 END i464
 PIN i465
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 189.72 174.70 190.28 ;
  END
 END i465
 PIN i466
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 185.53 174.70 186.10 ;
  END
 END i466
 PIN i467
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 181.54 174.70 182.12 ;
  END
 END i467
 PIN i468
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 177.37 174.70 177.94 ;
  END
 END i468
 PIN i469
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 778.34 174.70 778.90 ;
  END
 END i469
 PIN i470
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 173.38 174.70 173.94 ;
  END
 END i470
 PIN i471
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 169.19 174.70 169.76 ;
  END
 END i471
 PIN i472
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 165.21 174.70 165.78 ;
  END
 END i472
 PIN i473
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 161.03 174.70 161.59 ;
  END
 END i473
 PIN i474
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 157.03 174.70 157.60 ;
  END
 END i474
 PIN i475
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 152.85 174.70 153.43 ;
  END
 END i475
 PIN i476
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 148.87 174.70 149.44 ;
  END
 END i476
 PIN i477
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 144.69 174.70 145.25 ;
  END
 END i477
 PIN i478
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 140.69 174.70 141.26 ;
  END
 END i478
 PIN i479
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 136.51 174.70 137.09 ;
  END
 END i479
 PIN i480
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 774.15 174.70 774.73 ;
  END
 END i480
 PIN i481
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 132.53 174.70 133.09 ;
  END
 END i481
 PIN i482
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 128.34 174.70 128.91 ;
  END
 END i482
 PIN i483
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 124.36 174.70 124.92 ;
  END
 END i483
 PIN i484
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 120.17 174.70 120.75 ;
  END
 END i484
 PIN i485
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 116.19 174.70 116.75 ;
  END
 END i485
 PIN i486
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 112.00 174.70 112.58 ;
  END
 END i486
 PIN i487
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 89.78 174.70 90.34 ;
  END
 END i487
 PIN i488
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 85.59 174.70 86.17 ;
  END
 END i488
 PIN i489
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 81.61 174.70 82.17 ;
  END
 END i489
 PIN i490
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 77.42 174.70 78.00 ;
  END
 END i490
 PIN i491
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 770.16 174.70 770.74 ;
  END
 END i491
 PIN i492
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 73.44 174.70 74.00 ;
  END
 END i492
 PIN i493
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 69.25 174.70 69.83 ;
  END
 END i493
 PIN i494
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 65.27 174.70 65.83 ;
  END
 END i494
 PIN i495
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 61.09 174.70 61.66 ;
  END
 END i495
 PIN i496
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 57.09 174.70 57.66 ;
  END
 END i496
 PIN i497
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 52.91 174.70 53.48 ;
  END
 END i497
 PIN i498
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 48.92 174.70 49.49 ;
  END
 END i498
 PIN i499
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 44.74 174.70 45.31 ;
  END
 END i499
 PIN i500
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 40.76 174.70 41.33 ;
  END
 END i500
 PIN i501
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 36.58 174.70 37.15 ;
  END
 END i501
 PIN i502
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 765.99 174.70 766.55 ;
  END
 END i502
 PIN i503
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 32.59 174.70 33.16 ;
  END
 END i503
 PIN i504
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 28.41 174.70 28.98 ;
  END
 END i504
 PIN i505
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 24.41 174.70 24.98 ;
  END
 END i505
 PIN i506
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 20.23 174.70 20.80 ;
  END
 END i506
 PIN i507
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 16.25 174.70 16.82 ;
  END
 END i507
 PIN i508
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 12.06 174.70 12.63 ;
  END
 END i508
 PIN i509
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 8.07 174.70 8.64 ;
  END
 END i509
 PIN i510
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 3.90 174.70 4.46 ;
  END
 END i510
 PIN i511
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 762.00 174.70 762.57 ;
  END
 END i511
 PIN i512
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 757.82 174.70 758.38 ;
  END
 END i512
 PIN i513
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 827.36 174.70 827.92 ;
  END
 END i513
 PIN i514
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 753.83 174.70 754.39 ;
  END
 END i514
 PIN i515
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 749.64 174.70 750.22 ;
  END
 END i515
 PIN i516
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 745.65 174.70 746.23 ;
  END
 END i516
 PIN i517
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 723.24 174.70 723.80 ;
  END
 END i517
 PIN i518
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 719.25 174.70 719.82 ;
  END
 END i518
 PIN i519
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 715.07 174.70 715.63 ;
  END
 END i519
 PIN i520
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 711.08 174.70 711.64 ;
  END
 END i520
 PIN i521
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 706.89 174.70 707.47 ;
  END
 END i521
 PIN i522
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 702.90 174.70 703.48 ;
  END
 END i522
 PIN i523
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 698.73 174.70 699.29 ;
  END
 END i523
 PIN i524
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 823.17 174.70 823.75 ;
  END
 END i524
 PIN i525
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 694.74 174.70 695.30 ;
  END
 END i525
 PIN i526
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 690.55 174.70 691.12 ;
  END
 END i526
 PIN i527
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 686.57 174.70 687.13 ;
  END
 END i527
 PIN i528
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 682.38 174.70 682.96 ;
  END
 END i528
 PIN i529
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 678.39 174.70 678.97 ;
  END
 END i529
 PIN i530
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 674.22 174.70 674.78 ;
  END
 END i530
 PIN i531
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 670.23 174.70 670.79 ;
  END
 END i531
 PIN i532
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 666.04 174.70 666.62 ;
  END
 END i532
 PIN i533
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 662.05 174.70 662.62 ;
  END
 END i533
 PIN i534
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 657.88 174.70 658.45 ;
  END
 END i534
 PIN i535
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 819.18 174.70 819.75 ;
  END
 END i535
 PIN i536
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 653.88 174.70 654.46 ;
  END
 END i536
 PIN i537
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 649.71 174.70 650.27 ;
  END
 END i537
 PIN i538
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 645.72 174.70 646.28 ;
  END
 END i538
 PIN i539
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 641.53 174.70 642.11 ;
  END
 END i539
 PIN i540
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 637.54 174.70 638.12 ;
  END
 END i540
 PIN i541
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 633.37 174.70 633.93 ;
  END
 END i541
 PIN i542
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 624.25 174.70 624.82 ;
  END
 END i542
 PIN i543
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 620.07 174.70 620.63 ;
  END
 END i543
 PIN i544
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 616.08 174.70 616.64 ;
  END
 END i544
 PIN i545
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 611.89 174.70 612.47 ;
  END
 END i545
 PIN i546
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 815.00 174.70 815.58 ;
  END
 END i546
 PIN i547
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 607.90 174.70 608.48 ;
  END
 END i547
 PIN i548
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 603.73 174.70 604.29 ;
  END
 END i548
 PIN i549
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 599.74 174.70 600.30 ;
  END
 END i549
 PIN i550
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 595.55 174.70 596.12 ;
  END
 END i550
 PIN i551
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 591.57 174.70 592.13 ;
  END
 END i551
 PIN i552
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 587.38 174.70 587.96 ;
  END
 END i552
 PIN i553
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 583.39 174.70 583.97 ;
  END
 END i553
 PIN i554
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 579.22 174.70 579.78 ;
  END
 END i554
 PIN i555
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 575.23 174.70 575.79 ;
  END
 END i555
 PIN i556
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 571.04 174.70 571.62 ;
  END
 END i556
 PIN i557
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 811.01 174.70 811.59 ;
  END
 END i557
 PIN i558
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 567.05 174.70 567.62 ;
  END
 END i558
 PIN i559
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 562.88 174.70 563.45 ;
  END
 END i559
 PIN i560
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 558.88 174.70 559.46 ;
  END
 END i560
 PIN i561
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 554.71 174.70 555.27 ;
  END
 END i561
 PIN i562
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 550.72 174.70 551.28 ;
  END
 END i562
 PIN i563
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 546.53 174.70 547.11 ;
  END
 END i563
 PIN i564
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 542.54 174.70 543.12 ;
  END
 END i564
 PIN i565
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 538.37 174.70 538.93 ;
  END
 END i565
 PIN i566
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 516.13 174.70 516.71 ;
  END
 END i566
 PIN i567
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 511.95 174.70 512.52 ;
  END
 END i567
 PIN i568
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 806.84 174.70 807.40 ;
  END
 END i568
 PIN i569
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 507.96 174.70 508.54 ;
  END
 END i569
 PIN i570
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 503.79 174.70 504.36 ;
  END
 END i570
 PIN i571
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 499.80 174.70 500.37 ;
  END
 END i571
 PIN i572
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 495.62 174.70 496.19 ;
  END
 END i572
 PIN i573
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 491.62 174.70 492.19 ;
  END
 END i573
 PIN i574
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 487.44 174.70 488.01 ;
  END
 END i574
 PIN i575
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 483.45 174.70 484.02 ;
  END
 END i575
 PIN i576
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 479.27 174.70 479.85 ;
  END
 END i576
 PIN i577
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 475.29 174.70 475.86 ;
  END
 END i577
 PIN i578
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 471.11 174.70 471.68 ;
  END
 END i578
 PIN i579
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 802.85 174.70 803.41 ;
  END
 END i579
 PIN i580
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 467.12 174.70 467.69 ;
  END
 END i580
 PIN i581
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 462.94 174.70 463.50 ;
  END
 END i581
 PIN i582
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 458.94 174.70 459.51 ;
  END
 END i582
 PIN i583
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 454.76 174.70 455.33 ;
  END
 END i583
 PIN i584
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 450.77 174.70 451.35 ;
  END
 END i584
 PIN i585
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 446.60 174.70 447.17 ;
  END
 END i585
 PIN i586
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 442.61 174.70 443.18 ;
  END
 END i586
 PIN i587
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 438.43 174.70 439.00 ;
  END
 END i587
 PIN i588
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 434.44 174.70 435.00 ;
  END
 END i588
 PIN i589
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 430.25 174.70 430.82 ;
  END
 END i589
 PIN i590
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 798.66 174.70 799.24 ;
  END
 END i590
 PIN i591
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 401.00 174.70 401.56 ;
  END
 END i591
 PIN i592
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 396.81 174.70 397.38 ;
  END
 END i592
 PIN i593
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 392.82 174.70 393.39 ;
  END
 END i593
 PIN i594
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 388.64 174.70 389.21 ;
  END
 END i594
 PIN i595
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 384.65 174.70 385.23 ;
  END
 END i595
 PIN i596
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 380.48 174.70 381.05 ;
  END
 END i596
 PIN i597
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 376.49 174.70 377.06 ;
  END
 END i597
 PIN i598
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 372.31 174.70 372.88 ;
  END
 END i598
 PIN i599
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 368.31 174.70 368.88 ;
  END
 END i599
 PIN i600
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 174.13 364.13 174.70 364.70 ;
  END
 END i600
 PIN i601
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 197.69 427.98 198.26 428.55 ;
  END
 END i601
 PIN i602
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 196.55 427.98 197.12 428.55 ;
  END
 END i602
 PIN i603
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 195.03 427.98 195.60 428.55 ;
  END
 END i603
 PIN i604
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 193.13 427.98 193.70 428.55 ;
  END
 END i604
 PIN i605
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 192.00 427.98 192.56 428.55 ;
  END
 END i605
 PIN i606
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 197.69 414.68 198.26 415.25 ;
  END
 END i606
 PIN i607
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 196.55 414.68 197.12 415.25 ;
  END
 END i607
 PIN i608
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 195.03 414.68 195.60 415.25 ;
  END
 END i608
 PIN i609
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 193.13 414.68 193.70 415.25 ;
  END
 END i609
 PIN i610
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 192.00 414.68 192.56 415.25 ;
  END
 END i610
 OBS
  LAYER metal1 ;
   RECT 0.00 0.00 179.36 1.71 ;
   RECT 0.00 1.71 179.36 3.42 ;
   RECT 0.00 3.42 179.36 5.13 ;
   RECT 0.00 5.13 179.36 6.84 ;
   RECT 0.00 6.84 179.36 8.55 ;
   RECT 0.00 8.55 179.36 10.26 ;
   RECT 0.00 10.26 179.36 11.97 ;
   RECT 0.00 11.97 179.36 13.68 ;
   RECT 0.00 13.68 179.36 15.39 ;
   RECT 0.00 15.39 179.36 17.10 ;
   RECT 0.00 17.10 179.36 18.81 ;
   RECT 0.00 18.81 179.36 20.52 ;
   RECT 0.00 20.52 179.36 22.23 ;
   RECT 0.00 22.23 179.36 23.94 ;
   RECT 0.00 23.94 179.36 25.65 ;
   RECT 0.00 25.65 179.36 27.36 ;
   RECT 0.00 27.36 179.36 29.07 ;
   RECT 0.00 29.07 179.36 30.78 ;
   RECT 0.00 30.78 179.36 32.49 ;
   RECT 0.00 32.49 179.36 34.20 ;
   RECT 0.00 34.20 179.36 35.91 ;
   RECT 0.00 35.91 179.36 37.62 ;
   RECT 0.00 37.62 179.36 39.33 ;
   RECT 0.00 39.33 179.36 41.04 ;
   RECT 0.00 41.04 179.36 42.75 ;
   RECT 0.00 42.75 179.36 44.46 ;
   RECT 0.00 44.46 179.36 46.17 ;
   RECT 0.00 46.17 179.36 47.88 ;
   RECT 0.00 47.88 179.36 49.59 ;
   RECT 0.00 49.59 179.36 51.30 ;
   RECT 0.00 51.30 179.36 53.01 ;
   RECT 0.00 53.01 179.36 54.72 ;
   RECT 0.00 54.72 179.36 56.43 ;
   RECT 0.00 56.43 179.36 58.14 ;
   RECT 0.00 58.14 179.36 59.85 ;
   RECT 0.00 59.85 179.36 61.56 ;
   RECT 0.00 61.56 179.36 63.27 ;
   RECT 0.00 63.27 179.36 64.98 ;
   RECT 0.00 64.98 179.36 66.69 ;
   RECT 0.00 66.69 179.36 68.40 ;
   RECT 0.00 68.40 179.36 70.11 ;
   RECT 0.00 70.11 179.36 71.82 ;
   RECT 0.00 71.82 179.36 73.53 ;
   RECT 0.00 73.53 179.36 75.24 ;
   RECT 0.00 75.24 179.36 76.95 ;
   RECT 0.00 76.95 179.36 78.66 ;
   RECT 0.00 78.66 179.36 80.37 ;
   RECT 0.00 80.37 179.36 82.08 ;
   RECT 0.00 82.08 179.36 83.79 ;
   RECT 0.00 83.79 179.36 85.50 ;
   RECT 0.00 85.50 179.36 87.21 ;
   RECT 0.00 87.21 179.36 88.92 ;
   RECT 0.00 88.92 179.36 90.63 ;
   RECT 0.00 90.63 179.36 92.34 ;
   RECT 0.00 92.34 179.36 94.05 ;
   RECT 0.00 94.05 179.36 95.76 ;
   RECT 0.00 95.76 179.36 97.47 ;
   RECT 0.00 97.47 179.36 99.18 ;
   RECT 0.00 99.18 179.36 100.89 ;
   RECT 0.00 100.89 179.36 102.60 ;
   RECT 0.00 102.60 179.36 104.31 ;
   RECT 0.00 104.31 179.36 106.02 ;
   RECT 0.00 106.02 179.36 107.73 ;
   RECT 0.00 107.73 179.36 109.44 ;
   RECT 0.00 109.44 179.36 111.15 ;
   RECT 0.00 111.15 179.36 112.86 ;
   RECT 0.00 112.86 179.36 114.57 ;
   RECT 0.00 114.57 179.36 116.28 ;
   RECT 0.00 116.28 179.36 117.99 ;
   RECT 0.00 117.99 179.36 119.70 ;
   RECT 0.00 119.70 179.36 121.41 ;
   RECT 0.00 121.41 179.36 123.12 ;
   RECT 0.00 123.12 179.36 124.83 ;
   RECT 0.00 124.83 179.36 126.54 ;
   RECT 0.00 126.54 179.36 128.25 ;
   RECT 0.00 128.25 179.36 129.96 ;
   RECT 0.00 129.96 179.36 131.67 ;
   RECT 0.00 131.67 179.36 133.38 ;
   RECT 0.00 133.38 179.36 135.09 ;
   RECT 0.00 135.09 179.36 136.80 ;
   RECT 0.00 136.80 179.36 138.51 ;
   RECT 0.00 138.51 179.36 140.22 ;
   RECT 0.00 140.22 179.36 141.93 ;
   RECT 0.00 141.93 179.36 143.64 ;
   RECT 0.00 143.64 179.36 145.35 ;
   RECT 0.00 145.35 179.36 147.06 ;
   RECT 0.00 147.06 179.36 148.77 ;
   RECT 0.00 148.77 179.36 150.48 ;
   RECT 0.00 150.48 179.36 152.19 ;
   RECT 0.00 152.19 179.36 153.90 ;
   RECT 0.00 153.90 179.36 155.61 ;
   RECT 0.00 155.61 179.36 157.32 ;
   RECT 0.00 157.32 179.36 159.03 ;
   RECT 0.00 159.03 179.36 160.74 ;
   RECT 0.00 160.74 179.36 162.45 ;
   RECT 0.00 162.45 179.36 164.16 ;
   RECT 0.00 164.16 179.36 165.87 ;
   RECT 0.00 165.87 179.36 167.58 ;
   RECT 0.00 167.58 179.36 169.29 ;
   RECT 0.00 169.29 179.36 171.00 ;
   RECT 0.00 171.00 179.36 172.71 ;
   RECT 0.00 172.71 179.36 174.42 ;
   RECT 0.00 174.42 179.36 176.13 ;
   RECT 0.00 176.13 179.36 177.84 ;
   RECT 0.00 177.84 179.36 179.55 ;
   RECT 0.00 179.55 179.36 181.26 ;
   RECT 0.00 181.26 179.36 182.97 ;
   RECT 0.00 182.97 179.36 184.68 ;
   RECT 0.00 184.68 179.36 186.39 ;
   RECT 0.00 186.39 179.36 188.10 ;
   RECT 0.00 188.10 179.36 189.81 ;
   RECT 0.00 189.81 179.36 191.52 ;
   RECT 0.00 191.52 179.36 193.23 ;
   RECT 0.00 193.23 179.36 194.94 ;
   RECT 0.00 194.94 179.36 196.65 ;
   RECT 0.00 196.65 179.36 198.36 ;
   RECT 0.00 198.36 179.36 200.07 ;
   RECT 0.00 200.07 179.36 201.78 ;
   RECT 0.00 201.78 179.36 203.49 ;
   RECT 0.00 203.49 179.36 205.20 ;
   RECT 0.00 205.20 179.36 206.91 ;
   RECT 0.00 206.91 179.36 208.62 ;
   RECT 0.00 208.62 179.36 210.33 ;
   RECT 0.00 210.33 179.36 212.04 ;
   RECT 0.00 212.04 179.36 213.75 ;
   RECT 0.00 213.75 179.36 215.46 ;
   RECT 0.00 215.46 179.36 217.17 ;
   RECT 0.00 217.17 179.36 218.88 ;
   RECT 0.00 218.88 179.36 220.59 ;
   RECT 0.00 220.59 179.36 222.30 ;
   RECT 0.00 222.30 179.36 224.01 ;
   RECT 0.00 224.01 179.36 225.72 ;
   RECT 0.00 225.72 179.36 227.43 ;
   RECT 0.00 227.43 179.36 229.14 ;
   RECT 0.00 229.14 179.36 230.85 ;
   RECT 0.00 230.85 179.36 232.56 ;
   RECT 0.00 232.56 179.36 234.27 ;
   RECT 0.00 234.27 179.36 235.98 ;
   RECT 0.00 235.98 179.36 237.69 ;
   RECT 0.00 237.69 179.36 239.40 ;
   RECT 0.00 239.40 179.36 241.11 ;
   RECT 0.00 241.11 179.36 242.82 ;
   RECT 0.00 242.82 179.36 244.53 ;
   RECT 0.00 244.53 179.36 246.24 ;
   RECT 0.00 246.24 179.36 247.95 ;
   RECT 0.00 247.95 179.36 249.66 ;
   RECT 0.00 249.66 179.36 251.37 ;
   RECT 0.00 251.37 179.36 253.08 ;
   RECT 0.00 253.08 179.36 254.79 ;
   RECT 0.00 254.79 179.36 256.50 ;
   RECT 0.00 256.50 179.36 258.21 ;
   RECT 0.00 258.21 179.36 259.92 ;
   RECT 0.00 259.92 179.36 261.63 ;
   RECT 0.00 261.63 179.36 263.34 ;
   RECT 0.00 263.34 179.36 265.05 ;
   RECT 0.00 265.05 179.36 266.76 ;
   RECT 0.00 266.76 179.36 268.47 ;
   RECT 0.00 268.47 179.36 270.18 ;
   RECT 0.00 270.18 179.36 271.89 ;
   RECT 0.00 271.89 179.36 273.60 ;
   RECT 0.00 273.60 179.36 275.31 ;
   RECT 0.00 275.31 179.36 277.02 ;
   RECT 0.00 277.02 179.36 278.73 ;
   RECT 0.00 278.73 179.36 280.44 ;
   RECT 0.00 280.44 179.36 282.15 ;
   RECT 0.00 282.15 179.36 283.86 ;
   RECT 0.00 283.86 179.36 285.57 ;
   RECT 0.00 285.57 179.36 287.28 ;
   RECT 0.00 287.28 179.36 288.99 ;
   RECT 0.00 288.99 179.36 290.70 ;
   RECT 0.00 290.70 179.36 292.41 ;
   RECT 0.00 292.41 179.36 294.12 ;
   RECT 0.00 294.12 179.36 295.83 ;
   RECT 0.00 295.83 179.36 297.54 ;
   RECT 0.00 297.54 179.36 299.25 ;
   RECT 0.00 299.25 179.36 300.96 ;
   RECT 0.00 300.96 179.36 302.67 ;
   RECT 0.00 302.67 179.36 304.38 ;
   RECT 0.00 304.38 179.36 306.09 ;
   RECT 0.00 306.09 179.36 307.80 ;
   RECT 0.00 307.80 179.36 309.51 ;
   RECT 0.00 309.51 179.36 311.22 ;
   RECT 0.00 311.22 179.36 312.93 ;
   RECT 0.00 312.93 179.36 314.64 ;
   RECT 0.00 314.64 179.36 316.35 ;
   RECT 0.00 316.35 179.36 318.06 ;
   RECT 0.00 318.06 179.36 319.77 ;
   RECT 0.00 319.77 179.36 321.48 ;
   RECT 0.00 321.48 179.36 323.19 ;
   RECT 0.00 323.19 179.36 324.90 ;
   RECT 0.00 324.90 179.36 326.61 ;
   RECT 0.00 326.61 179.36 328.32 ;
   RECT 0.00 328.32 179.36 330.03 ;
   RECT 0.00 330.03 179.36 331.74 ;
   RECT 0.00 331.74 179.36 333.45 ;
   RECT 0.00 333.45 179.36 335.16 ;
   RECT 0.00 335.16 179.36 336.87 ;
   RECT 0.00 336.87 179.36 338.58 ;
   RECT 0.00 338.58 179.36 340.29 ;
   RECT 0.00 340.29 179.36 342.00 ;
   RECT 0.00 342.00 179.36 343.71 ;
   RECT 0.00 343.71 179.36 345.42 ;
   RECT 0.00 345.42 179.36 347.13 ;
   RECT 0.00 347.13 179.36 348.84 ;
   RECT 0.00 348.84 179.36 350.55 ;
   RECT 0.00 350.55 179.36 352.26 ;
   RECT 0.00 352.26 179.36 353.97 ;
   RECT 0.00 353.97 179.36 355.68 ;
   RECT 0.00 355.68 179.36 357.39 ;
   RECT 0.00 357.39 179.36 359.10 ;
   RECT 0.00 359.10 179.36 360.81 ;
   RECT 0.00 360.81 179.36 362.52 ;
   RECT 0.00 362.52 179.36 364.23 ;
   RECT 0.00 364.23 179.36 365.94 ;
   RECT 0.00 365.94 179.36 367.65 ;
   RECT 0.00 367.65 179.36 369.36 ;
   RECT 0.00 369.36 179.36 371.07 ;
   RECT 0.00 371.07 179.36 372.78 ;
   RECT 0.00 372.78 179.36 374.49 ;
   RECT 0.00 374.49 179.36 376.20 ;
   RECT 0.00 376.20 179.36 377.91 ;
   RECT 0.00 377.91 179.36 379.62 ;
   RECT 0.00 379.62 179.36 381.33 ;
   RECT 0.00 381.33 179.36 383.04 ;
   RECT 0.00 383.04 179.36 384.75 ;
   RECT 0.00 384.75 179.36 386.46 ;
   RECT 0.00 386.46 179.36 388.17 ;
   RECT 0.00 388.17 179.36 389.88 ;
   RECT 0.00 389.88 179.36 391.59 ;
   RECT 0.00 391.59 179.36 393.30 ;
   RECT 0.00 393.30 179.36 395.01 ;
   RECT 0.00 395.01 179.36 396.72 ;
   RECT 0.00 396.72 179.36 398.43 ;
   RECT 0.00 398.43 179.36 400.14 ;
   RECT 0.00 400.14 179.36 401.85 ;
   RECT 0.00 401.85 202.54 403.56 ;
   RECT 0.00 403.56 202.54 405.27 ;
   RECT 0.00 405.27 202.54 406.98 ;
   RECT 0.00 406.98 202.54 408.69 ;
   RECT 0.00 408.69 202.54 410.40 ;
   RECT 0.00 410.40 202.54 412.11 ;
   RECT 0.00 412.11 202.54 413.82 ;
   RECT 0.00 413.82 202.54 415.53 ;
   RECT 0.00 415.53 202.54 417.24 ;
   RECT 0.00 417.24 202.54 418.95 ;
   RECT 0.00 418.95 202.54 420.66 ;
   RECT 0.00 420.66 202.54 422.37 ;
   RECT 0.00 422.37 202.54 424.08 ;
   RECT 0.00 424.08 202.54 425.79 ;
   RECT 0.00 425.79 202.54 427.50 ;
   RECT 0.00 427.50 202.54 429.21 ;
   RECT 0.00 429.21 202.54 430.92 ;
   RECT 0.00 430.92 179.36 432.63 ;
   RECT 0.00 432.63 179.36 434.34 ;
   RECT 0.00 434.34 179.36 436.05 ;
   RECT 0.00 436.05 179.36 437.76 ;
   RECT 0.00 437.76 179.36 439.47 ;
   RECT 0.00 439.47 179.36 441.18 ;
   RECT 0.00 441.18 179.36 442.89 ;
   RECT 0.00 442.89 179.36 444.60 ;
   RECT 0.00 444.60 179.36 446.31 ;
   RECT 0.00 446.31 179.36 448.02 ;
   RECT 0.00 448.02 179.36 449.73 ;
   RECT 0.00 449.73 179.36 451.44 ;
   RECT 0.00 451.44 179.36 453.15 ;
   RECT 0.00 453.15 179.36 454.86 ;
   RECT 0.00 454.86 179.36 456.57 ;
   RECT 0.00 456.57 179.36 458.28 ;
   RECT 0.00 458.28 179.36 459.99 ;
   RECT 0.00 459.99 179.36 461.70 ;
   RECT 0.00 461.70 179.36 463.41 ;
   RECT 0.00 463.41 179.36 465.12 ;
   RECT 0.00 465.12 179.36 466.83 ;
   RECT 0.00 466.83 179.36 468.54 ;
   RECT 0.00 468.54 179.36 470.25 ;
   RECT 0.00 470.25 179.36 471.96 ;
   RECT 0.00 471.96 179.36 473.67 ;
   RECT 0.00 473.67 179.36 475.38 ;
   RECT 0.00 475.38 179.36 477.09 ;
   RECT 0.00 477.09 179.36 478.80 ;
   RECT 0.00 478.80 179.36 480.51 ;
   RECT 0.00 480.51 179.36 482.22 ;
   RECT 0.00 482.22 179.36 483.93 ;
   RECT 0.00 483.93 179.36 485.64 ;
   RECT 0.00 485.64 179.36 487.35 ;
   RECT 0.00 487.35 179.36 489.06 ;
   RECT 0.00 489.06 179.36 490.77 ;
   RECT 0.00 490.77 179.36 492.48 ;
   RECT 0.00 492.48 179.36 494.19 ;
   RECT 0.00 494.19 179.36 495.90 ;
   RECT 0.00 495.90 179.36 497.61 ;
   RECT 0.00 497.61 179.36 499.32 ;
   RECT 0.00 499.32 179.36 501.03 ;
   RECT 0.00 501.03 179.36 502.74 ;
   RECT 0.00 502.74 179.36 504.45 ;
   RECT 0.00 504.45 179.36 506.16 ;
   RECT 0.00 506.16 179.36 507.87 ;
   RECT 0.00 507.87 179.36 509.58 ;
   RECT 0.00 509.58 179.36 511.29 ;
   RECT 0.00 511.29 179.36 513.00 ;
   RECT 0.00 513.00 179.36 514.71 ;
   RECT 0.00 514.71 179.36 516.42 ;
   RECT 0.00 516.42 179.36 518.13 ;
   RECT 0.00 518.13 179.36 519.84 ;
   RECT 0.00 519.84 179.36 521.55 ;
   RECT 0.00 521.55 179.36 523.26 ;
   RECT 0.00 523.26 179.36 524.97 ;
   RECT 0.00 524.97 179.36 526.68 ;
   RECT 0.00 526.68 179.36 528.39 ;
   RECT 0.00 528.39 179.36 530.10 ;
   RECT 0.00 530.10 179.36 531.81 ;
   RECT 0.00 531.81 179.36 533.52 ;
   RECT 0.00 533.52 179.36 535.23 ;
   RECT 0.00 535.23 179.36 536.94 ;
   RECT 0.00 536.94 179.36 538.65 ;
   RECT 0.00 538.65 179.36 540.36 ;
   RECT 0.00 540.36 179.36 542.07 ;
   RECT 0.00 542.07 179.36 543.78 ;
   RECT 0.00 543.78 179.36 545.49 ;
   RECT 0.00 545.49 179.36 547.20 ;
   RECT 0.00 547.20 179.36 548.91 ;
   RECT 0.00 548.91 179.36 550.62 ;
   RECT 0.00 550.62 179.36 552.33 ;
   RECT 0.00 552.33 179.36 554.04 ;
   RECT 0.00 554.04 179.36 555.75 ;
   RECT 0.00 555.75 179.36 557.46 ;
   RECT 0.00 557.46 179.36 559.17 ;
   RECT 0.00 559.17 179.36 560.88 ;
   RECT 0.00 560.88 179.36 562.59 ;
   RECT 0.00 562.59 179.36 564.30 ;
   RECT 0.00 564.30 179.36 566.01 ;
   RECT 0.00 566.01 179.36 567.72 ;
   RECT 0.00 567.72 179.36 569.43 ;
   RECT 0.00 569.43 179.36 571.14 ;
   RECT 0.00 571.14 179.36 572.85 ;
   RECT 0.00 572.85 179.36 574.56 ;
   RECT 0.00 574.56 179.36 576.27 ;
   RECT 0.00 576.27 179.36 577.98 ;
   RECT 0.00 577.98 179.36 579.69 ;
   RECT 0.00 579.69 179.36 581.40 ;
   RECT 0.00 581.40 179.36 583.11 ;
   RECT 0.00 583.11 179.36 584.82 ;
   RECT 0.00 584.82 179.36 586.53 ;
   RECT 0.00 586.53 179.36 588.24 ;
   RECT 0.00 588.24 179.36 589.95 ;
   RECT 0.00 589.95 179.36 591.66 ;
   RECT 0.00 591.66 179.36 593.37 ;
   RECT 0.00 593.37 179.36 595.08 ;
   RECT 0.00 595.08 179.36 596.79 ;
   RECT 0.00 596.79 179.36 598.50 ;
   RECT 0.00 598.50 179.36 600.21 ;
   RECT 0.00 600.21 179.36 601.92 ;
   RECT 0.00 601.92 179.36 603.63 ;
   RECT 0.00 603.63 179.36 605.34 ;
   RECT 0.00 605.34 179.36 607.05 ;
   RECT 0.00 607.05 179.36 608.76 ;
   RECT 0.00 608.76 179.36 610.47 ;
   RECT 0.00 610.47 179.36 612.18 ;
   RECT 0.00 612.18 179.36 613.89 ;
   RECT 0.00 613.89 179.36 615.60 ;
   RECT 0.00 615.60 179.36 617.31 ;
   RECT 0.00 617.31 179.36 619.02 ;
   RECT 0.00 619.02 179.36 620.73 ;
   RECT 0.00 620.73 179.36 622.44 ;
   RECT 0.00 622.44 179.36 624.15 ;
   RECT 0.00 624.15 179.36 625.86 ;
   RECT 0.00 625.86 179.36 627.57 ;
   RECT 0.00 627.57 179.36 629.28 ;
   RECT 0.00 629.28 179.36 630.99 ;
   RECT 0.00 630.99 179.36 632.70 ;
   RECT 0.00 632.70 179.36 634.41 ;
   RECT 0.00 634.41 179.36 636.12 ;
   RECT 0.00 636.12 179.36 637.83 ;
   RECT 0.00 637.83 179.36 639.54 ;
   RECT 0.00 639.54 179.36 641.25 ;
   RECT 0.00 641.25 179.36 642.96 ;
   RECT 0.00 642.96 179.36 644.67 ;
   RECT 0.00 644.67 179.36 646.38 ;
   RECT 0.00 646.38 179.36 648.09 ;
   RECT 0.00 648.09 179.36 649.80 ;
   RECT 0.00 649.80 179.36 651.51 ;
   RECT 0.00 651.51 179.36 653.22 ;
   RECT 0.00 653.22 179.36 654.93 ;
   RECT 0.00 654.93 179.36 656.64 ;
   RECT 0.00 656.64 179.36 658.35 ;
   RECT 0.00 658.35 179.36 660.06 ;
   RECT 0.00 660.06 179.36 661.77 ;
   RECT 0.00 661.77 179.36 663.48 ;
   RECT 0.00 663.48 179.36 665.19 ;
   RECT 0.00 665.19 179.36 666.90 ;
   RECT 0.00 666.90 179.36 668.61 ;
   RECT 0.00 668.61 179.36 670.32 ;
   RECT 0.00 670.32 179.36 672.03 ;
   RECT 0.00 672.03 179.36 673.74 ;
   RECT 0.00 673.74 179.36 675.45 ;
   RECT 0.00 675.45 179.36 677.16 ;
   RECT 0.00 677.16 179.36 678.87 ;
   RECT 0.00 678.87 179.36 680.58 ;
   RECT 0.00 680.58 179.36 682.29 ;
   RECT 0.00 682.29 179.36 684.00 ;
   RECT 0.00 684.00 179.36 685.71 ;
   RECT 0.00 685.71 179.36 687.42 ;
   RECT 0.00 687.42 179.36 689.13 ;
   RECT 0.00 689.13 179.36 690.84 ;
   RECT 0.00 690.84 179.36 692.55 ;
   RECT 0.00 692.55 179.36 694.26 ;
   RECT 0.00 694.26 179.36 695.97 ;
   RECT 0.00 695.97 179.36 697.68 ;
   RECT 0.00 697.68 179.36 699.39 ;
   RECT 0.00 699.39 179.36 701.10 ;
   RECT 0.00 701.10 179.36 702.81 ;
   RECT 0.00 702.81 179.36 704.52 ;
   RECT 0.00 704.52 179.36 706.23 ;
   RECT 0.00 706.23 179.36 707.94 ;
   RECT 0.00 707.94 179.36 709.65 ;
   RECT 0.00 709.65 179.36 711.36 ;
   RECT 0.00 711.36 179.36 713.07 ;
   RECT 0.00 713.07 179.36 714.78 ;
   RECT 0.00 714.78 179.36 716.49 ;
   RECT 0.00 716.49 179.36 718.20 ;
   RECT 0.00 718.20 179.36 719.91 ;
   RECT 0.00 719.91 179.36 721.62 ;
   RECT 0.00 721.62 179.36 723.33 ;
   RECT 0.00 723.33 179.36 725.04 ;
   RECT 0.00 725.04 179.36 726.75 ;
   RECT 0.00 726.75 179.36 728.46 ;
   RECT 0.00 728.46 179.36 730.17 ;
   RECT 0.00 730.17 179.36 731.88 ;
   RECT 0.00 731.88 179.36 733.59 ;
   RECT 0.00 733.59 179.36 735.30 ;
   RECT 0.00 735.30 179.36 737.01 ;
   RECT 0.00 737.01 179.36 738.72 ;
   RECT 0.00 738.72 179.36 740.43 ;
   RECT 0.00 740.43 179.36 742.14 ;
   RECT 0.00 742.14 179.36 743.85 ;
   RECT 0.00 743.85 179.36 745.56 ;
   RECT 0.00 745.56 179.36 747.27 ;
   RECT 0.00 747.27 179.36 748.98 ;
   RECT 0.00 748.98 179.36 750.69 ;
   RECT 0.00 750.69 179.36 752.40 ;
   RECT 0.00 752.40 179.36 754.11 ;
   RECT 0.00 754.11 179.36 755.82 ;
   RECT 0.00 755.82 179.36 757.53 ;
   RECT 0.00 757.53 179.36 759.24 ;
   RECT 0.00 759.24 179.36 760.95 ;
   RECT 0.00 760.95 179.36 762.66 ;
   RECT 0.00 762.66 179.36 764.37 ;
   RECT 0.00 764.37 179.36 766.08 ;
   RECT 0.00 766.08 179.36 767.79 ;
   RECT 0.00 767.79 179.36 769.50 ;
   RECT 0.00 769.50 179.36 771.21 ;
   RECT 0.00 771.21 179.36 772.92 ;
   RECT 0.00 772.92 179.36 774.63 ;
   RECT 0.00 774.63 179.36 776.34 ;
   RECT 0.00 776.34 179.36 778.05 ;
   RECT 0.00 778.05 179.36 779.76 ;
   RECT 0.00 779.76 179.36 781.47 ;
   RECT 0.00 781.47 179.36 783.18 ;
   RECT 0.00 783.18 179.36 784.89 ;
   RECT 0.00 784.89 179.36 786.60 ;
   RECT 0.00 786.60 179.36 788.31 ;
   RECT 0.00 788.31 179.36 790.02 ;
   RECT 0.00 790.02 179.36 791.73 ;
   RECT 0.00 791.73 179.36 793.44 ;
   RECT 0.00 793.44 179.36 795.15 ;
   RECT 0.00 795.15 179.36 796.86 ;
   RECT 0.00 796.86 179.36 798.57 ;
   RECT 0.00 798.57 179.36 800.28 ;
   RECT 0.00 800.28 179.36 801.99 ;
   RECT 0.00 801.99 179.36 803.70 ;
   RECT 0.00 803.70 179.36 805.41 ;
   RECT 0.00 805.41 179.36 807.12 ;
   RECT 0.00 807.12 179.36 808.83 ;
   RECT 0.00 808.83 179.36 810.54 ;
   RECT 0.00 810.54 179.36 812.25 ;
   RECT 0.00 812.25 179.36 813.96 ;
   RECT 0.00 813.96 179.36 815.67 ;
   RECT 0.00 815.67 179.36 817.38 ;
   RECT 0.00 817.38 179.36 819.09 ;
   RECT 0.00 819.09 179.36 820.80 ;
   RECT 0.00 820.80 179.36 822.51 ;
   RECT 0.00 822.51 179.36 824.22 ;
   RECT 0.00 824.22 179.36 825.93 ;
   RECT 0.00 825.93 179.36 827.64 ;
   RECT 0.00 827.64 179.36 829.35 ;
   RECT 0.00 829.35 179.36 831.06 ;
   RECT 0.00 831.06 179.36 832.77 ;
   RECT 0.00 832.77 179.36 834.48 ;
   RECT 0.00 834.48 179.36 836.19 ;
   RECT 0.00 836.19 179.36 837.90 ;
   RECT 0.00 837.90 179.36 839.61 ;
   RECT 0.00 839.61 179.36 841.32 ;
  LAYER via1 ;
   RECT 0.00 0.00 179.36 1.71 ;
   RECT 0.00 1.71 179.36 3.42 ;
   RECT 0.00 3.42 179.36 5.13 ;
   RECT 0.00 5.13 179.36 6.84 ;
   RECT 0.00 6.84 179.36 8.55 ;
   RECT 0.00 8.55 179.36 10.26 ;
   RECT 0.00 10.26 179.36 11.97 ;
   RECT 0.00 11.97 179.36 13.68 ;
   RECT 0.00 13.68 179.36 15.39 ;
   RECT 0.00 15.39 179.36 17.10 ;
   RECT 0.00 17.10 179.36 18.81 ;
   RECT 0.00 18.81 179.36 20.52 ;
   RECT 0.00 20.52 179.36 22.23 ;
   RECT 0.00 22.23 179.36 23.94 ;
   RECT 0.00 23.94 179.36 25.65 ;
   RECT 0.00 25.65 179.36 27.36 ;
   RECT 0.00 27.36 179.36 29.07 ;
   RECT 0.00 29.07 179.36 30.78 ;
   RECT 0.00 30.78 179.36 32.49 ;
   RECT 0.00 32.49 179.36 34.20 ;
   RECT 0.00 34.20 179.36 35.91 ;
   RECT 0.00 35.91 179.36 37.62 ;
   RECT 0.00 37.62 179.36 39.33 ;
   RECT 0.00 39.33 179.36 41.04 ;
   RECT 0.00 41.04 179.36 42.75 ;
   RECT 0.00 42.75 179.36 44.46 ;
   RECT 0.00 44.46 179.36 46.17 ;
   RECT 0.00 46.17 179.36 47.88 ;
   RECT 0.00 47.88 179.36 49.59 ;
   RECT 0.00 49.59 179.36 51.30 ;
   RECT 0.00 51.30 179.36 53.01 ;
   RECT 0.00 53.01 179.36 54.72 ;
   RECT 0.00 54.72 179.36 56.43 ;
   RECT 0.00 56.43 179.36 58.14 ;
   RECT 0.00 58.14 179.36 59.85 ;
   RECT 0.00 59.85 179.36 61.56 ;
   RECT 0.00 61.56 179.36 63.27 ;
   RECT 0.00 63.27 179.36 64.98 ;
   RECT 0.00 64.98 179.36 66.69 ;
   RECT 0.00 66.69 179.36 68.40 ;
   RECT 0.00 68.40 179.36 70.11 ;
   RECT 0.00 70.11 179.36 71.82 ;
   RECT 0.00 71.82 179.36 73.53 ;
   RECT 0.00 73.53 179.36 75.24 ;
   RECT 0.00 75.24 179.36 76.95 ;
   RECT 0.00 76.95 179.36 78.66 ;
   RECT 0.00 78.66 179.36 80.37 ;
   RECT 0.00 80.37 179.36 82.08 ;
   RECT 0.00 82.08 179.36 83.79 ;
   RECT 0.00 83.79 179.36 85.50 ;
   RECT 0.00 85.50 179.36 87.21 ;
   RECT 0.00 87.21 179.36 88.92 ;
   RECT 0.00 88.92 179.36 90.63 ;
   RECT 0.00 90.63 179.36 92.34 ;
   RECT 0.00 92.34 179.36 94.05 ;
   RECT 0.00 94.05 179.36 95.76 ;
   RECT 0.00 95.76 179.36 97.47 ;
   RECT 0.00 97.47 179.36 99.18 ;
   RECT 0.00 99.18 179.36 100.89 ;
   RECT 0.00 100.89 179.36 102.60 ;
   RECT 0.00 102.60 179.36 104.31 ;
   RECT 0.00 104.31 179.36 106.02 ;
   RECT 0.00 106.02 179.36 107.73 ;
   RECT 0.00 107.73 179.36 109.44 ;
   RECT 0.00 109.44 179.36 111.15 ;
   RECT 0.00 111.15 179.36 112.86 ;
   RECT 0.00 112.86 179.36 114.57 ;
   RECT 0.00 114.57 179.36 116.28 ;
   RECT 0.00 116.28 179.36 117.99 ;
   RECT 0.00 117.99 179.36 119.70 ;
   RECT 0.00 119.70 179.36 121.41 ;
   RECT 0.00 121.41 179.36 123.12 ;
   RECT 0.00 123.12 179.36 124.83 ;
   RECT 0.00 124.83 179.36 126.54 ;
   RECT 0.00 126.54 179.36 128.25 ;
   RECT 0.00 128.25 179.36 129.96 ;
   RECT 0.00 129.96 179.36 131.67 ;
   RECT 0.00 131.67 179.36 133.38 ;
   RECT 0.00 133.38 179.36 135.09 ;
   RECT 0.00 135.09 179.36 136.80 ;
   RECT 0.00 136.80 179.36 138.51 ;
   RECT 0.00 138.51 179.36 140.22 ;
   RECT 0.00 140.22 179.36 141.93 ;
   RECT 0.00 141.93 179.36 143.64 ;
   RECT 0.00 143.64 179.36 145.35 ;
   RECT 0.00 145.35 179.36 147.06 ;
   RECT 0.00 147.06 179.36 148.77 ;
   RECT 0.00 148.77 179.36 150.48 ;
   RECT 0.00 150.48 179.36 152.19 ;
   RECT 0.00 152.19 179.36 153.90 ;
   RECT 0.00 153.90 179.36 155.61 ;
   RECT 0.00 155.61 179.36 157.32 ;
   RECT 0.00 157.32 179.36 159.03 ;
   RECT 0.00 159.03 179.36 160.74 ;
   RECT 0.00 160.74 179.36 162.45 ;
   RECT 0.00 162.45 179.36 164.16 ;
   RECT 0.00 164.16 179.36 165.87 ;
   RECT 0.00 165.87 179.36 167.58 ;
   RECT 0.00 167.58 179.36 169.29 ;
   RECT 0.00 169.29 179.36 171.00 ;
   RECT 0.00 171.00 179.36 172.71 ;
   RECT 0.00 172.71 179.36 174.42 ;
   RECT 0.00 174.42 179.36 176.13 ;
   RECT 0.00 176.13 179.36 177.84 ;
   RECT 0.00 177.84 179.36 179.55 ;
   RECT 0.00 179.55 179.36 181.26 ;
   RECT 0.00 181.26 179.36 182.97 ;
   RECT 0.00 182.97 179.36 184.68 ;
   RECT 0.00 184.68 179.36 186.39 ;
   RECT 0.00 186.39 179.36 188.10 ;
   RECT 0.00 188.10 179.36 189.81 ;
   RECT 0.00 189.81 179.36 191.52 ;
   RECT 0.00 191.52 179.36 193.23 ;
   RECT 0.00 193.23 179.36 194.94 ;
   RECT 0.00 194.94 179.36 196.65 ;
   RECT 0.00 196.65 179.36 198.36 ;
   RECT 0.00 198.36 179.36 200.07 ;
   RECT 0.00 200.07 179.36 201.78 ;
   RECT 0.00 201.78 179.36 203.49 ;
   RECT 0.00 203.49 179.36 205.20 ;
   RECT 0.00 205.20 179.36 206.91 ;
   RECT 0.00 206.91 179.36 208.62 ;
   RECT 0.00 208.62 179.36 210.33 ;
   RECT 0.00 210.33 179.36 212.04 ;
   RECT 0.00 212.04 179.36 213.75 ;
   RECT 0.00 213.75 179.36 215.46 ;
   RECT 0.00 215.46 179.36 217.17 ;
   RECT 0.00 217.17 179.36 218.88 ;
   RECT 0.00 218.88 179.36 220.59 ;
   RECT 0.00 220.59 179.36 222.30 ;
   RECT 0.00 222.30 179.36 224.01 ;
   RECT 0.00 224.01 179.36 225.72 ;
   RECT 0.00 225.72 179.36 227.43 ;
   RECT 0.00 227.43 179.36 229.14 ;
   RECT 0.00 229.14 179.36 230.85 ;
   RECT 0.00 230.85 179.36 232.56 ;
   RECT 0.00 232.56 179.36 234.27 ;
   RECT 0.00 234.27 179.36 235.98 ;
   RECT 0.00 235.98 179.36 237.69 ;
   RECT 0.00 237.69 179.36 239.40 ;
   RECT 0.00 239.40 179.36 241.11 ;
   RECT 0.00 241.11 179.36 242.82 ;
   RECT 0.00 242.82 179.36 244.53 ;
   RECT 0.00 244.53 179.36 246.24 ;
   RECT 0.00 246.24 179.36 247.95 ;
   RECT 0.00 247.95 179.36 249.66 ;
   RECT 0.00 249.66 179.36 251.37 ;
   RECT 0.00 251.37 179.36 253.08 ;
   RECT 0.00 253.08 179.36 254.79 ;
   RECT 0.00 254.79 179.36 256.50 ;
   RECT 0.00 256.50 179.36 258.21 ;
   RECT 0.00 258.21 179.36 259.92 ;
   RECT 0.00 259.92 179.36 261.63 ;
   RECT 0.00 261.63 179.36 263.34 ;
   RECT 0.00 263.34 179.36 265.05 ;
   RECT 0.00 265.05 179.36 266.76 ;
   RECT 0.00 266.76 179.36 268.47 ;
   RECT 0.00 268.47 179.36 270.18 ;
   RECT 0.00 270.18 179.36 271.89 ;
   RECT 0.00 271.89 179.36 273.60 ;
   RECT 0.00 273.60 179.36 275.31 ;
   RECT 0.00 275.31 179.36 277.02 ;
   RECT 0.00 277.02 179.36 278.73 ;
   RECT 0.00 278.73 179.36 280.44 ;
   RECT 0.00 280.44 179.36 282.15 ;
   RECT 0.00 282.15 179.36 283.86 ;
   RECT 0.00 283.86 179.36 285.57 ;
   RECT 0.00 285.57 179.36 287.28 ;
   RECT 0.00 287.28 179.36 288.99 ;
   RECT 0.00 288.99 179.36 290.70 ;
   RECT 0.00 290.70 179.36 292.41 ;
   RECT 0.00 292.41 179.36 294.12 ;
   RECT 0.00 294.12 179.36 295.83 ;
   RECT 0.00 295.83 179.36 297.54 ;
   RECT 0.00 297.54 179.36 299.25 ;
   RECT 0.00 299.25 179.36 300.96 ;
   RECT 0.00 300.96 179.36 302.67 ;
   RECT 0.00 302.67 179.36 304.38 ;
   RECT 0.00 304.38 179.36 306.09 ;
   RECT 0.00 306.09 179.36 307.80 ;
   RECT 0.00 307.80 179.36 309.51 ;
   RECT 0.00 309.51 179.36 311.22 ;
   RECT 0.00 311.22 179.36 312.93 ;
   RECT 0.00 312.93 179.36 314.64 ;
   RECT 0.00 314.64 179.36 316.35 ;
   RECT 0.00 316.35 179.36 318.06 ;
   RECT 0.00 318.06 179.36 319.77 ;
   RECT 0.00 319.77 179.36 321.48 ;
   RECT 0.00 321.48 179.36 323.19 ;
   RECT 0.00 323.19 179.36 324.90 ;
   RECT 0.00 324.90 179.36 326.61 ;
   RECT 0.00 326.61 179.36 328.32 ;
   RECT 0.00 328.32 179.36 330.03 ;
   RECT 0.00 330.03 179.36 331.74 ;
   RECT 0.00 331.74 179.36 333.45 ;
   RECT 0.00 333.45 179.36 335.16 ;
   RECT 0.00 335.16 179.36 336.87 ;
   RECT 0.00 336.87 179.36 338.58 ;
   RECT 0.00 338.58 179.36 340.29 ;
   RECT 0.00 340.29 179.36 342.00 ;
   RECT 0.00 342.00 179.36 343.71 ;
   RECT 0.00 343.71 179.36 345.42 ;
   RECT 0.00 345.42 179.36 347.13 ;
   RECT 0.00 347.13 179.36 348.84 ;
   RECT 0.00 348.84 179.36 350.55 ;
   RECT 0.00 350.55 179.36 352.26 ;
   RECT 0.00 352.26 179.36 353.97 ;
   RECT 0.00 353.97 179.36 355.68 ;
   RECT 0.00 355.68 179.36 357.39 ;
   RECT 0.00 357.39 179.36 359.10 ;
   RECT 0.00 359.10 179.36 360.81 ;
   RECT 0.00 360.81 179.36 362.52 ;
   RECT 0.00 362.52 179.36 364.23 ;
   RECT 0.00 364.23 179.36 365.94 ;
   RECT 0.00 365.94 179.36 367.65 ;
   RECT 0.00 367.65 179.36 369.36 ;
   RECT 0.00 369.36 179.36 371.07 ;
   RECT 0.00 371.07 179.36 372.78 ;
   RECT 0.00 372.78 179.36 374.49 ;
   RECT 0.00 374.49 179.36 376.20 ;
   RECT 0.00 376.20 179.36 377.91 ;
   RECT 0.00 377.91 179.36 379.62 ;
   RECT 0.00 379.62 179.36 381.33 ;
   RECT 0.00 381.33 179.36 383.04 ;
   RECT 0.00 383.04 179.36 384.75 ;
   RECT 0.00 384.75 179.36 386.46 ;
   RECT 0.00 386.46 179.36 388.17 ;
   RECT 0.00 388.17 179.36 389.88 ;
   RECT 0.00 389.88 179.36 391.59 ;
   RECT 0.00 391.59 179.36 393.30 ;
   RECT 0.00 393.30 179.36 395.01 ;
   RECT 0.00 395.01 179.36 396.72 ;
   RECT 0.00 396.72 179.36 398.43 ;
   RECT 0.00 398.43 179.36 400.14 ;
   RECT 0.00 400.14 179.36 401.85 ;
   RECT 0.00 401.85 202.54 403.56 ;
   RECT 0.00 403.56 202.54 405.27 ;
   RECT 0.00 405.27 202.54 406.98 ;
   RECT 0.00 406.98 202.54 408.69 ;
   RECT 0.00 408.69 202.54 410.40 ;
   RECT 0.00 410.40 202.54 412.11 ;
   RECT 0.00 412.11 202.54 413.82 ;
   RECT 0.00 413.82 202.54 415.53 ;
   RECT 0.00 415.53 202.54 417.24 ;
   RECT 0.00 417.24 202.54 418.95 ;
   RECT 0.00 418.95 202.54 420.66 ;
   RECT 0.00 420.66 202.54 422.37 ;
   RECT 0.00 422.37 202.54 424.08 ;
   RECT 0.00 424.08 202.54 425.79 ;
   RECT 0.00 425.79 202.54 427.50 ;
   RECT 0.00 427.50 202.54 429.21 ;
   RECT 0.00 429.21 202.54 430.92 ;
   RECT 0.00 430.92 179.36 432.63 ;
   RECT 0.00 432.63 179.36 434.34 ;
   RECT 0.00 434.34 179.36 436.05 ;
   RECT 0.00 436.05 179.36 437.76 ;
   RECT 0.00 437.76 179.36 439.47 ;
   RECT 0.00 439.47 179.36 441.18 ;
   RECT 0.00 441.18 179.36 442.89 ;
   RECT 0.00 442.89 179.36 444.60 ;
   RECT 0.00 444.60 179.36 446.31 ;
   RECT 0.00 446.31 179.36 448.02 ;
   RECT 0.00 448.02 179.36 449.73 ;
   RECT 0.00 449.73 179.36 451.44 ;
   RECT 0.00 451.44 179.36 453.15 ;
   RECT 0.00 453.15 179.36 454.86 ;
   RECT 0.00 454.86 179.36 456.57 ;
   RECT 0.00 456.57 179.36 458.28 ;
   RECT 0.00 458.28 179.36 459.99 ;
   RECT 0.00 459.99 179.36 461.70 ;
   RECT 0.00 461.70 179.36 463.41 ;
   RECT 0.00 463.41 179.36 465.12 ;
   RECT 0.00 465.12 179.36 466.83 ;
   RECT 0.00 466.83 179.36 468.54 ;
   RECT 0.00 468.54 179.36 470.25 ;
   RECT 0.00 470.25 179.36 471.96 ;
   RECT 0.00 471.96 179.36 473.67 ;
   RECT 0.00 473.67 179.36 475.38 ;
   RECT 0.00 475.38 179.36 477.09 ;
   RECT 0.00 477.09 179.36 478.80 ;
   RECT 0.00 478.80 179.36 480.51 ;
   RECT 0.00 480.51 179.36 482.22 ;
   RECT 0.00 482.22 179.36 483.93 ;
   RECT 0.00 483.93 179.36 485.64 ;
   RECT 0.00 485.64 179.36 487.35 ;
   RECT 0.00 487.35 179.36 489.06 ;
   RECT 0.00 489.06 179.36 490.77 ;
   RECT 0.00 490.77 179.36 492.48 ;
   RECT 0.00 492.48 179.36 494.19 ;
   RECT 0.00 494.19 179.36 495.90 ;
   RECT 0.00 495.90 179.36 497.61 ;
   RECT 0.00 497.61 179.36 499.32 ;
   RECT 0.00 499.32 179.36 501.03 ;
   RECT 0.00 501.03 179.36 502.74 ;
   RECT 0.00 502.74 179.36 504.45 ;
   RECT 0.00 504.45 179.36 506.16 ;
   RECT 0.00 506.16 179.36 507.87 ;
   RECT 0.00 507.87 179.36 509.58 ;
   RECT 0.00 509.58 179.36 511.29 ;
   RECT 0.00 511.29 179.36 513.00 ;
   RECT 0.00 513.00 179.36 514.71 ;
   RECT 0.00 514.71 179.36 516.42 ;
   RECT 0.00 516.42 179.36 518.13 ;
   RECT 0.00 518.13 179.36 519.84 ;
   RECT 0.00 519.84 179.36 521.55 ;
   RECT 0.00 521.55 179.36 523.26 ;
   RECT 0.00 523.26 179.36 524.97 ;
   RECT 0.00 524.97 179.36 526.68 ;
   RECT 0.00 526.68 179.36 528.39 ;
   RECT 0.00 528.39 179.36 530.10 ;
   RECT 0.00 530.10 179.36 531.81 ;
   RECT 0.00 531.81 179.36 533.52 ;
   RECT 0.00 533.52 179.36 535.23 ;
   RECT 0.00 535.23 179.36 536.94 ;
   RECT 0.00 536.94 179.36 538.65 ;
   RECT 0.00 538.65 179.36 540.36 ;
   RECT 0.00 540.36 179.36 542.07 ;
   RECT 0.00 542.07 179.36 543.78 ;
   RECT 0.00 543.78 179.36 545.49 ;
   RECT 0.00 545.49 179.36 547.20 ;
   RECT 0.00 547.20 179.36 548.91 ;
   RECT 0.00 548.91 179.36 550.62 ;
   RECT 0.00 550.62 179.36 552.33 ;
   RECT 0.00 552.33 179.36 554.04 ;
   RECT 0.00 554.04 179.36 555.75 ;
   RECT 0.00 555.75 179.36 557.46 ;
   RECT 0.00 557.46 179.36 559.17 ;
   RECT 0.00 559.17 179.36 560.88 ;
   RECT 0.00 560.88 179.36 562.59 ;
   RECT 0.00 562.59 179.36 564.30 ;
   RECT 0.00 564.30 179.36 566.01 ;
   RECT 0.00 566.01 179.36 567.72 ;
   RECT 0.00 567.72 179.36 569.43 ;
   RECT 0.00 569.43 179.36 571.14 ;
   RECT 0.00 571.14 179.36 572.85 ;
   RECT 0.00 572.85 179.36 574.56 ;
   RECT 0.00 574.56 179.36 576.27 ;
   RECT 0.00 576.27 179.36 577.98 ;
   RECT 0.00 577.98 179.36 579.69 ;
   RECT 0.00 579.69 179.36 581.40 ;
   RECT 0.00 581.40 179.36 583.11 ;
   RECT 0.00 583.11 179.36 584.82 ;
   RECT 0.00 584.82 179.36 586.53 ;
   RECT 0.00 586.53 179.36 588.24 ;
   RECT 0.00 588.24 179.36 589.95 ;
   RECT 0.00 589.95 179.36 591.66 ;
   RECT 0.00 591.66 179.36 593.37 ;
   RECT 0.00 593.37 179.36 595.08 ;
   RECT 0.00 595.08 179.36 596.79 ;
   RECT 0.00 596.79 179.36 598.50 ;
   RECT 0.00 598.50 179.36 600.21 ;
   RECT 0.00 600.21 179.36 601.92 ;
   RECT 0.00 601.92 179.36 603.63 ;
   RECT 0.00 603.63 179.36 605.34 ;
   RECT 0.00 605.34 179.36 607.05 ;
   RECT 0.00 607.05 179.36 608.76 ;
   RECT 0.00 608.76 179.36 610.47 ;
   RECT 0.00 610.47 179.36 612.18 ;
   RECT 0.00 612.18 179.36 613.89 ;
   RECT 0.00 613.89 179.36 615.60 ;
   RECT 0.00 615.60 179.36 617.31 ;
   RECT 0.00 617.31 179.36 619.02 ;
   RECT 0.00 619.02 179.36 620.73 ;
   RECT 0.00 620.73 179.36 622.44 ;
   RECT 0.00 622.44 179.36 624.15 ;
   RECT 0.00 624.15 179.36 625.86 ;
   RECT 0.00 625.86 179.36 627.57 ;
   RECT 0.00 627.57 179.36 629.28 ;
   RECT 0.00 629.28 179.36 630.99 ;
   RECT 0.00 630.99 179.36 632.70 ;
   RECT 0.00 632.70 179.36 634.41 ;
   RECT 0.00 634.41 179.36 636.12 ;
   RECT 0.00 636.12 179.36 637.83 ;
   RECT 0.00 637.83 179.36 639.54 ;
   RECT 0.00 639.54 179.36 641.25 ;
   RECT 0.00 641.25 179.36 642.96 ;
   RECT 0.00 642.96 179.36 644.67 ;
   RECT 0.00 644.67 179.36 646.38 ;
   RECT 0.00 646.38 179.36 648.09 ;
   RECT 0.00 648.09 179.36 649.80 ;
   RECT 0.00 649.80 179.36 651.51 ;
   RECT 0.00 651.51 179.36 653.22 ;
   RECT 0.00 653.22 179.36 654.93 ;
   RECT 0.00 654.93 179.36 656.64 ;
   RECT 0.00 656.64 179.36 658.35 ;
   RECT 0.00 658.35 179.36 660.06 ;
   RECT 0.00 660.06 179.36 661.77 ;
   RECT 0.00 661.77 179.36 663.48 ;
   RECT 0.00 663.48 179.36 665.19 ;
   RECT 0.00 665.19 179.36 666.90 ;
   RECT 0.00 666.90 179.36 668.61 ;
   RECT 0.00 668.61 179.36 670.32 ;
   RECT 0.00 670.32 179.36 672.03 ;
   RECT 0.00 672.03 179.36 673.74 ;
   RECT 0.00 673.74 179.36 675.45 ;
   RECT 0.00 675.45 179.36 677.16 ;
   RECT 0.00 677.16 179.36 678.87 ;
   RECT 0.00 678.87 179.36 680.58 ;
   RECT 0.00 680.58 179.36 682.29 ;
   RECT 0.00 682.29 179.36 684.00 ;
   RECT 0.00 684.00 179.36 685.71 ;
   RECT 0.00 685.71 179.36 687.42 ;
   RECT 0.00 687.42 179.36 689.13 ;
   RECT 0.00 689.13 179.36 690.84 ;
   RECT 0.00 690.84 179.36 692.55 ;
   RECT 0.00 692.55 179.36 694.26 ;
   RECT 0.00 694.26 179.36 695.97 ;
   RECT 0.00 695.97 179.36 697.68 ;
   RECT 0.00 697.68 179.36 699.39 ;
   RECT 0.00 699.39 179.36 701.10 ;
   RECT 0.00 701.10 179.36 702.81 ;
   RECT 0.00 702.81 179.36 704.52 ;
   RECT 0.00 704.52 179.36 706.23 ;
   RECT 0.00 706.23 179.36 707.94 ;
   RECT 0.00 707.94 179.36 709.65 ;
   RECT 0.00 709.65 179.36 711.36 ;
   RECT 0.00 711.36 179.36 713.07 ;
   RECT 0.00 713.07 179.36 714.78 ;
   RECT 0.00 714.78 179.36 716.49 ;
   RECT 0.00 716.49 179.36 718.20 ;
   RECT 0.00 718.20 179.36 719.91 ;
   RECT 0.00 719.91 179.36 721.62 ;
   RECT 0.00 721.62 179.36 723.33 ;
   RECT 0.00 723.33 179.36 725.04 ;
   RECT 0.00 725.04 179.36 726.75 ;
   RECT 0.00 726.75 179.36 728.46 ;
   RECT 0.00 728.46 179.36 730.17 ;
   RECT 0.00 730.17 179.36 731.88 ;
   RECT 0.00 731.88 179.36 733.59 ;
   RECT 0.00 733.59 179.36 735.30 ;
   RECT 0.00 735.30 179.36 737.01 ;
   RECT 0.00 737.01 179.36 738.72 ;
   RECT 0.00 738.72 179.36 740.43 ;
   RECT 0.00 740.43 179.36 742.14 ;
   RECT 0.00 742.14 179.36 743.85 ;
   RECT 0.00 743.85 179.36 745.56 ;
   RECT 0.00 745.56 179.36 747.27 ;
   RECT 0.00 747.27 179.36 748.98 ;
   RECT 0.00 748.98 179.36 750.69 ;
   RECT 0.00 750.69 179.36 752.40 ;
   RECT 0.00 752.40 179.36 754.11 ;
   RECT 0.00 754.11 179.36 755.82 ;
   RECT 0.00 755.82 179.36 757.53 ;
   RECT 0.00 757.53 179.36 759.24 ;
   RECT 0.00 759.24 179.36 760.95 ;
   RECT 0.00 760.95 179.36 762.66 ;
   RECT 0.00 762.66 179.36 764.37 ;
   RECT 0.00 764.37 179.36 766.08 ;
   RECT 0.00 766.08 179.36 767.79 ;
   RECT 0.00 767.79 179.36 769.50 ;
   RECT 0.00 769.50 179.36 771.21 ;
   RECT 0.00 771.21 179.36 772.92 ;
   RECT 0.00 772.92 179.36 774.63 ;
   RECT 0.00 774.63 179.36 776.34 ;
   RECT 0.00 776.34 179.36 778.05 ;
   RECT 0.00 778.05 179.36 779.76 ;
   RECT 0.00 779.76 179.36 781.47 ;
   RECT 0.00 781.47 179.36 783.18 ;
   RECT 0.00 783.18 179.36 784.89 ;
   RECT 0.00 784.89 179.36 786.60 ;
   RECT 0.00 786.60 179.36 788.31 ;
   RECT 0.00 788.31 179.36 790.02 ;
   RECT 0.00 790.02 179.36 791.73 ;
   RECT 0.00 791.73 179.36 793.44 ;
   RECT 0.00 793.44 179.36 795.15 ;
   RECT 0.00 795.15 179.36 796.86 ;
   RECT 0.00 796.86 179.36 798.57 ;
   RECT 0.00 798.57 179.36 800.28 ;
   RECT 0.00 800.28 179.36 801.99 ;
   RECT 0.00 801.99 179.36 803.70 ;
   RECT 0.00 803.70 179.36 805.41 ;
   RECT 0.00 805.41 179.36 807.12 ;
   RECT 0.00 807.12 179.36 808.83 ;
   RECT 0.00 808.83 179.36 810.54 ;
   RECT 0.00 810.54 179.36 812.25 ;
   RECT 0.00 812.25 179.36 813.96 ;
   RECT 0.00 813.96 179.36 815.67 ;
   RECT 0.00 815.67 179.36 817.38 ;
   RECT 0.00 817.38 179.36 819.09 ;
   RECT 0.00 819.09 179.36 820.80 ;
   RECT 0.00 820.80 179.36 822.51 ;
   RECT 0.00 822.51 179.36 824.22 ;
   RECT 0.00 824.22 179.36 825.93 ;
   RECT 0.00 825.93 179.36 827.64 ;
   RECT 0.00 827.64 179.36 829.35 ;
   RECT 0.00 829.35 179.36 831.06 ;
   RECT 0.00 831.06 179.36 832.77 ;
   RECT 0.00 832.77 179.36 834.48 ;
   RECT 0.00 834.48 179.36 836.19 ;
   RECT 0.00 836.19 179.36 837.90 ;
   RECT 0.00 837.90 179.36 839.61 ;
   RECT 0.00 839.61 179.36 841.32 ;
  LAYER metal2 ;
   RECT 0.00 0.00 179.36 1.71 ;
   RECT 0.00 1.71 179.36 3.42 ;
   RECT 0.00 3.42 179.36 5.13 ;
   RECT 0.00 5.13 179.36 6.84 ;
   RECT 0.00 6.84 179.36 8.55 ;
   RECT 0.00 8.55 179.36 10.26 ;
   RECT 0.00 10.26 179.36 11.97 ;
   RECT 0.00 11.97 179.36 13.68 ;
   RECT 0.00 13.68 179.36 15.39 ;
   RECT 0.00 15.39 179.36 17.10 ;
   RECT 0.00 17.10 179.36 18.81 ;
   RECT 0.00 18.81 179.36 20.52 ;
   RECT 0.00 20.52 179.36 22.23 ;
   RECT 0.00 22.23 179.36 23.94 ;
   RECT 0.00 23.94 179.36 25.65 ;
   RECT 0.00 25.65 179.36 27.36 ;
   RECT 0.00 27.36 179.36 29.07 ;
   RECT 0.00 29.07 179.36 30.78 ;
   RECT 0.00 30.78 179.36 32.49 ;
   RECT 0.00 32.49 179.36 34.20 ;
   RECT 0.00 34.20 179.36 35.91 ;
   RECT 0.00 35.91 179.36 37.62 ;
   RECT 0.00 37.62 179.36 39.33 ;
   RECT 0.00 39.33 179.36 41.04 ;
   RECT 0.00 41.04 179.36 42.75 ;
   RECT 0.00 42.75 179.36 44.46 ;
   RECT 0.00 44.46 179.36 46.17 ;
   RECT 0.00 46.17 179.36 47.88 ;
   RECT 0.00 47.88 179.36 49.59 ;
   RECT 0.00 49.59 179.36 51.30 ;
   RECT 0.00 51.30 179.36 53.01 ;
   RECT 0.00 53.01 179.36 54.72 ;
   RECT 0.00 54.72 179.36 56.43 ;
   RECT 0.00 56.43 179.36 58.14 ;
   RECT 0.00 58.14 179.36 59.85 ;
   RECT 0.00 59.85 179.36 61.56 ;
   RECT 0.00 61.56 179.36 63.27 ;
   RECT 0.00 63.27 179.36 64.98 ;
   RECT 0.00 64.98 179.36 66.69 ;
   RECT 0.00 66.69 179.36 68.40 ;
   RECT 0.00 68.40 179.36 70.11 ;
   RECT 0.00 70.11 179.36 71.82 ;
   RECT 0.00 71.82 179.36 73.53 ;
   RECT 0.00 73.53 179.36 75.24 ;
   RECT 0.00 75.24 179.36 76.95 ;
   RECT 0.00 76.95 179.36 78.66 ;
   RECT 0.00 78.66 179.36 80.37 ;
   RECT 0.00 80.37 179.36 82.08 ;
   RECT 0.00 82.08 179.36 83.79 ;
   RECT 0.00 83.79 179.36 85.50 ;
   RECT 0.00 85.50 179.36 87.21 ;
   RECT 0.00 87.21 179.36 88.92 ;
   RECT 0.00 88.92 179.36 90.63 ;
   RECT 0.00 90.63 179.36 92.34 ;
   RECT 0.00 92.34 179.36 94.05 ;
   RECT 0.00 94.05 179.36 95.76 ;
   RECT 0.00 95.76 179.36 97.47 ;
   RECT 0.00 97.47 179.36 99.18 ;
   RECT 0.00 99.18 179.36 100.89 ;
   RECT 0.00 100.89 179.36 102.60 ;
   RECT 0.00 102.60 179.36 104.31 ;
   RECT 0.00 104.31 179.36 106.02 ;
   RECT 0.00 106.02 179.36 107.73 ;
   RECT 0.00 107.73 179.36 109.44 ;
   RECT 0.00 109.44 179.36 111.15 ;
   RECT 0.00 111.15 179.36 112.86 ;
   RECT 0.00 112.86 179.36 114.57 ;
   RECT 0.00 114.57 179.36 116.28 ;
   RECT 0.00 116.28 179.36 117.99 ;
   RECT 0.00 117.99 179.36 119.70 ;
   RECT 0.00 119.70 179.36 121.41 ;
   RECT 0.00 121.41 179.36 123.12 ;
   RECT 0.00 123.12 179.36 124.83 ;
   RECT 0.00 124.83 179.36 126.54 ;
   RECT 0.00 126.54 179.36 128.25 ;
   RECT 0.00 128.25 179.36 129.96 ;
   RECT 0.00 129.96 179.36 131.67 ;
   RECT 0.00 131.67 179.36 133.38 ;
   RECT 0.00 133.38 179.36 135.09 ;
   RECT 0.00 135.09 179.36 136.80 ;
   RECT 0.00 136.80 179.36 138.51 ;
   RECT 0.00 138.51 179.36 140.22 ;
   RECT 0.00 140.22 179.36 141.93 ;
   RECT 0.00 141.93 179.36 143.64 ;
   RECT 0.00 143.64 179.36 145.35 ;
   RECT 0.00 145.35 179.36 147.06 ;
   RECT 0.00 147.06 179.36 148.77 ;
   RECT 0.00 148.77 179.36 150.48 ;
   RECT 0.00 150.48 179.36 152.19 ;
   RECT 0.00 152.19 179.36 153.90 ;
   RECT 0.00 153.90 179.36 155.61 ;
   RECT 0.00 155.61 179.36 157.32 ;
   RECT 0.00 157.32 179.36 159.03 ;
   RECT 0.00 159.03 179.36 160.74 ;
   RECT 0.00 160.74 179.36 162.45 ;
   RECT 0.00 162.45 179.36 164.16 ;
   RECT 0.00 164.16 179.36 165.87 ;
   RECT 0.00 165.87 179.36 167.58 ;
   RECT 0.00 167.58 179.36 169.29 ;
   RECT 0.00 169.29 179.36 171.00 ;
   RECT 0.00 171.00 179.36 172.71 ;
   RECT 0.00 172.71 179.36 174.42 ;
   RECT 0.00 174.42 179.36 176.13 ;
   RECT 0.00 176.13 179.36 177.84 ;
   RECT 0.00 177.84 179.36 179.55 ;
   RECT 0.00 179.55 179.36 181.26 ;
   RECT 0.00 181.26 179.36 182.97 ;
   RECT 0.00 182.97 179.36 184.68 ;
   RECT 0.00 184.68 179.36 186.39 ;
   RECT 0.00 186.39 179.36 188.10 ;
   RECT 0.00 188.10 179.36 189.81 ;
   RECT 0.00 189.81 179.36 191.52 ;
   RECT 0.00 191.52 179.36 193.23 ;
   RECT 0.00 193.23 179.36 194.94 ;
   RECT 0.00 194.94 179.36 196.65 ;
   RECT 0.00 196.65 179.36 198.36 ;
   RECT 0.00 198.36 179.36 200.07 ;
   RECT 0.00 200.07 179.36 201.78 ;
   RECT 0.00 201.78 179.36 203.49 ;
   RECT 0.00 203.49 179.36 205.20 ;
   RECT 0.00 205.20 179.36 206.91 ;
   RECT 0.00 206.91 179.36 208.62 ;
   RECT 0.00 208.62 179.36 210.33 ;
   RECT 0.00 210.33 179.36 212.04 ;
   RECT 0.00 212.04 179.36 213.75 ;
   RECT 0.00 213.75 179.36 215.46 ;
   RECT 0.00 215.46 179.36 217.17 ;
   RECT 0.00 217.17 179.36 218.88 ;
   RECT 0.00 218.88 179.36 220.59 ;
   RECT 0.00 220.59 179.36 222.30 ;
   RECT 0.00 222.30 179.36 224.01 ;
   RECT 0.00 224.01 179.36 225.72 ;
   RECT 0.00 225.72 179.36 227.43 ;
   RECT 0.00 227.43 179.36 229.14 ;
   RECT 0.00 229.14 179.36 230.85 ;
   RECT 0.00 230.85 179.36 232.56 ;
   RECT 0.00 232.56 179.36 234.27 ;
   RECT 0.00 234.27 179.36 235.98 ;
   RECT 0.00 235.98 179.36 237.69 ;
   RECT 0.00 237.69 179.36 239.40 ;
   RECT 0.00 239.40 179.36 241.11 ;
   RECT 0.00 241.11 179.36 242.82 ;
   RECT 0.00 242.82 179.36 244.53 ;
   RECT 0.00 244.53 179.36 246.24 ;
   RECT 0.00 246.24 179.36 247.95 ;
   RECT 0.00 247.95 179.36 249.66 ;
   RECT 0.00 249.66 179.36 251.37 ;
   RECT 0.00 251.37 179.36 253.08 ;
   RECT 0.00 253.08 179.36 254.79 ;
   RECT 0.00 254.79 179.36 256.50 ;
   RECT 0.00 256.50 179.36 258.21 ;
   RECT 0.00 258.21 179.36 259.92 ;
   RECT 0.00 259.92 179.36 261.63 ;
   RECT 0.00 261.63 179.36 263.34 ;
   RECT 0.00 263.34 179.36 265.05 ;
   RECT 0.00 265.05 179.36 266.76 ;
   RECT 0.00 266.76 179.36 268.47 ;
   RECT 0.00 268.47 179.36 270.18 ;
   RECT 0.00 270.18 179.36 271.89 ;
   RECT 0.00 271.89 179.36 273.60 ;
   RECT 0.00 273.60 179.36 275.31 ;
   RECT 0.00 275.31 179.36 277.02 ;
   RECT 0.00 277.02 179.36 278.73 ;
   RECT 0.00 278.73 179.36 280.44 ;
   RECT 0.00 280.44 179.36 282.15 ;
   RECT 0.00 282.15 179.36 283.86 ;
   RECT 0.00 283.86 179.36 285.57 ;
   RECT 0.00 285.57 179.36 287.28 ;
   RECT 0.00 287.28 179.36 288.99 ;
   RECT 0.00 288.99 179.36 290.70 ;
   RECT 0.00 290.70 179.36 292.41 ;
   RECT 0.00 292.41 179.36 294.12 ;
   RECT 0.00 294.12 179.36 295.83 ;
   RECT 0.00 295.83 179.36 297.54 ;
   RECT 0.00 297.54 179.36 299.25 ;
   RECT 0.00 299.25 179.36 300.96 ;
   RECT 0.00 300.96 179.36 302.67 ;
   RECT 0.00 302.67 179.36 304.38 ;
   RECT 0.00 304.38 179.36 306.09 ;
   RECT 0.00 306.09 179.36 307.80 ;
   RECT 0.00 307.80 179.36 309.51 ;
   RECT 0.00 309.51 179.36 311.22 ;
   RECT 0.00 311.22 179.36 312.93 ;
   RECT 0.00 312.93 179.36 314.64 ;
   RECT 0.00 314.64 179.36 316.35 ;
   RECT 0.00 316.35 179.36 318.06 ;
   RECT 0.00 318.06 179.36 319.77 ;
   RECT 0.00 319.77 179.36 321.48 ;
   RECT 0.00 321.48 179.36 323.19 ;
   RECT 0.00 323.19 179.36 324.90 ;
   RECT 0.00 324.90 179.36 326.61 ;
   RECT 0.00 326.61 179.36 328.32 ;
   RECT 0.00 328.32 179.36 330.03 ;
   RECT 0.00 330.03 179.36 331.74 ;
   RECT 0.00 331.74 179.36 333.45 ;
   RECT 0.00 333.45 179.36 335.16 ;
   RECT 0.00 335.16 179.36 336.87 ;
   RECT 0.00 336.87 179.36 338.58 ;
   RECT 0.00 338.58 179.36 340.29 ;
   RECT 0.00 340.29 179.36 342.00 ;
   RECT 0.00 342.00 179.36 343.71 ;
   RECT 0.00 343.71 179.36 345.42 ;
   RECT 0.00 345.42 179.36 347.13 ;
   RECT 0.00 347.13 179.36 348.84 ;
   RECT 0.00 348.84 179.36 350.55 ;
   RECT 0.00 350.55 179.36 352.26 ;
   RECT 0.00 352.26 179.36 353.97 ;
   RECT 0.00 353.97 179.36 355.68 ;
   RECT 0.00 355.68 179.36 357.39 ;
   RECT 0.00 357.39 179.36 359.10 ;
   RECT 0.00 359.10 179.36 360.81 ;
   RECT 0.00 360.81 179.36 362.52 ;
   RECT 0.00 362.52 179.36 364.23 ;
   RECT 0.00 364.23 179.36 365.94 ;
   RECT 0.00 365.94 179.36 367.65 ;
   RECT 0.00 367.65 179.36 369.36 ;
   RECT 0.00 369.36 179.36 371.07 ;
   RECT 0.00 371.07 179.36 372.78 ;
   RECT 0.00 372.78 179.36 374.49 ;
   RECT 0.00 374.49 179.36 376.20 ;
   RECT 0.00 376.20 179.36 377.91 ;
   RECT 0.00 377.91 179.36 379.62 ;
   RECT 0.00 379.62 179.36 381.33 ;
   RECT 0.00 381.33 179.36 383.04 ;
   RECT 0.00 383.04 179.36 384.75 ;
   RECT 0.00 384.75 179.36 386.46 ;
   RECT 0.00 386.46 179.36 388.17 ;
   RECT 0.00 388.17 179.36 389.88 ;
   RECT 0.00 389.88 179.36 391.59 ;
   RECT 0.00 391.59 179.36 393.30 ;
   RECT 0.00 393.30 179.36 395.01 ;
   RECT 0.00 395.01 179.36 396.72 ;
   RECT 0.00 396.72 179.36 398.43 ;
   RECT 0.00 398.43 179.36 400.14 ;
   RECT 0.00 400.14 179.36 401.85 ;
   RECT 0.00 401.85 202.54 403.56 ;
   RECT 0.00 403.56 202.54 405.27 ;
   RECT 0.00 405.27 202.54 406.98 ;
   RECT 0.00 406.98 202.54 408.69 ;
   RECT 0.00 408.69 202.54 410.40 ;
   RECT 0.00 410.40 202.54 412.11 ;
   RECT 0.00 412.11 202.54 413.82 ;
   RECT 0.00 413.82 202.54 415.53 ;
   RECT 0.00 415.53 202.54 417.24 ;
   RECT 0.00 417.24 202.54 418.95 ;
   RECT 0.00 418.95 202.54 420.66 ;
   RECT 0.00 420.66 202.54 422.37 ;
   RECT 0.00 422.37 202.54 424.08 ;
   RECT 0.00 424.08 202.54 425.79 ;
   RECT 0.00 425.79 202.54 427.50 ;
   RECT 0.00 427.50 202.54 429.21 ;
   RECT 0.00 429.21 202.54 430.92 ;
   RECT 0.00 430.92 179.36 432.63 ;
   RECT 0.00 432.63 179.36 434.34 ;
   RECT 0.00 434.34 179.36 436.05 ;
   RECT 0.00 436.05 179.36 437.76 ;
   RECT 0.00 437.76 179.36 439.47 ;
   RECT 0.00 439.47 179.36 441.18 ;
   RECT 0.00 441.18 179.36 442.89 ;
   RECT 0.00 442.89 179.36 444.60 ;
   RECT 0.00 444.60 179.36 446.31 ;
   RECT 0.00 446.31 179.36 448.02 ;
   RECT 0.00 448.02 179.36 449.73 ;
   RECT 0.00 449.73 179.36 451.44 ;
   RECT 0.00 451.44 179.36 453.15 ;
   RECT 0.00 453.15 179.36 454.86 ;
   RECT 0.00 454.86 179.36 456.57 ;
   RECT 0.00 456.57 179.36 458.28 ;
   RECT 0.00 458.28 179.36 459.99 ;
   RECT 0.00 459.99 179.36 461.70 ;
   RECT 0.00 461.70 179.36 463.41 ;
   RECT 0.00 463.41 179.36 465.12 ;
   RECT 0.00 465.12 179.36 466.83 ;
   RECT 0.00 466.83 179.36 468.54 ;
   RECT 0.00 468.54 179.36 470.25 ;
   RECT 0.00 470.25 179.36 471.96 ;
   RECT 0.00 471.96 179.36 473.67 ;
   RECT 0.00 473.67 179.36 475.38 ;
   RECT 0.00 475.38 179.36 477.09 ;
   RECT 0.00 477.09 179.36 478.80 ;
   RECT 0.00 478.80 179.36 480.51 ;
   RECT 0.00 480.51 179.36 482.22 ;
   RECT 0.00 482.22 179.36 483.93 ;
   RECT 0.00 483.93 179.36 485.64 ;
   RECT 0.00 485.64 179.36 487.35 ;
   RECT 0.00 487.35 179.36 489.06 ;
   RECT 0.00 489.06 179.36 490.77 ;
   RECT 0.00 490.77 179.36 492.48 ;
   RECT 0.00 492.48 179.36 494.19 ;
   RECT 0.00 494.19 179.36 495.90 ;
   RECT 0.00 495.90 179.36 497.61 ;
   RECT 0.00 497.61 179.36 499.32 ;
   RECT 0.00 499.32 179.36 501.03 ;
   RECT 0.00 501.03 179.36 502.74 ;
   RECT 0.00 502.74 179.36 504.45 ;
   RECT 0.00 504.45 179.36 506.16 ;
   RECT 0.00 506.16 179.36 507.87 ;
   RECT 0.00 507.87 179.36 509.58 ;
   RECT 0.00 509.58 179.36 511.29 ;
   RECT 0.00 511.29 179.36 513.00 ;
   RECT 0.00 513.00 179.36 514.71 ;
   RECT 0.00 514.71 179.36 516.42 ;
   RECT 0.00 516.42 179.36 518.13 ;
   RECT 0.00 518.13 179.36 519.84 ;
   RECT 0.00 519.84 179.36 521.55 ;
   RECT 0.00 521.55 179.36 523.26 ;
   RECT 0.00 523.26 179.36 524.97 ;
   RECT 0.00 524.97 179.36 526.68 ;
   RECT 0.00 526.68 179.36 528.39 ;
   RECT 0.00 528.39 179.36 530.10 ;
   RECT 0.00 530.10 179.36 531.81 ;
   RECT 0.00 531.81 179.36 533.52 ;
   RECT 0.00 533.52 179.36 535.23 ;
   RECT 0.00 535.23 179.36 536.94 ;
   RECT 0.00 536.94 179.36 538.65 ;
   RECT 0.00 538.65 179.36 540.36 ;
   RECT 0.00 540.36 179.36 542.07 ;
   RECT 0.00 542.07 179.36 543.78 ;
   RECT 0.00 543.78 179.36 545.49 ;
   RECT 0.00 545.49 179.36 547.20 ;
   RECT 0.00 547.20 179.36 548.91 ;
   RECT 0.00 548.91 179.36 550.62 ;
   RECT 0.00 550.62 179.36 552.33 ;
   RECT 0.00 552.33 179.36 554.04 ;
   RECT 0.00 554.04 179.36 555.75 ;
   RECT 0.00 555.75 179.36 557.46 ;
   RECT 0.00 557.46 179.36 559.17 ;
   RECT 0.00 559.17 179.36 560.88 ;
   RECT 0.00 560.88 179.36 562.59 ;
   RECT 0.00 562.59 179.36 564.30 ;
   RECT 0.00 564.30 179.36 566.01 ;
   RECT 0.00 566.01 179.36 567.72 ;
   RECT 0.00 567.72 179.36 569.43 ;
   RECT 0.00 569.43 179.36 571.14 ;
   RECT 0.00 571.14 179.36 572.85 ;
   RECT 0.00 572.85 179.36 574.56 ;
   RECT 0.00 574.56 179.36 576.27 ;
   RECT 0.00 576.27 179.36 577.98 ;
   RECT 0.00 577.98 179.36 579.69 ;
   RECT 0.00 579.69 179.36 581.40 ;
   RECT 0.00 581.40 179.36 583.11 ;
   RECT 0.00 583.11 179.36 584.82 ;
   RECT 0.00 584.82 179.36 586.53 ;
   RECT 0.00 586.53 179.36 588.24 ;
   RECT 0.00 588.24 179.36 589.95 ;
   RECT 0.00 589.95 179.36 591.66 ;
   RECT 0.00 591.66 179.36 593.37 ;
   RECT 0.00 593.37 179.36 595.08 ;
   RECT 0.00 595.08 179.36 596.79 ;
   RECT 0.00 596.79 179.36 598.50 ;
   RECT 0.00 598.50 179.36 600.21 ;
   RECT 0.00 600.21 179.36 601.92 ;
   RECT 0.00 601.92 179.36 603.63 ;
   RECT 0.00 603.63 179.36 605.34 ;
   RECT 0.00 605.34 179.36 607.05 ;
   RECT 0.00 607.05 179.36 608.76 ;
   RECT 0.00 608.76 179.36 610.47 ;
   RECT 0.00 610.47 179.36 612.18 ;
   RECT 0.00 612.18 179.36 613.89 ;
   RECT 0.00 613.89 179.36 615.60 ;
   RECT 0.00 615.60 179.36 617.31 ;
   RECT 0.00 617.31 179.36 619.02 ;
   RECT 0.00 619.02 179.36 620.73 ;
   RECT 0.00 620.73 179.36 622.44 ;
   RECT 0.00 622.44 179.36 624.15 ;
   RECT 0.00 624.15 179.36 625.86 ;
   RECT 0.00 625.86 179.36 627.57 ;
   RECT 0.00 627.57 179.36 629.28 ;
   RECT 0.00 629.28 179.36 630.99 ;
   RECT 0.00 630.99 179.36 632.70 ;
   RECT 0.00 632.70 179.36 634.41 ;
   RECT 0.00 634.41 179.36 636.12 ;
   RECT 0.00 636.12 179.36 637.83 ;
   RECT 0.00 637.83 179.36 639.54 ;
   RECT 0.00 639.54 179.36 641.25 ;
   RECT 0.00 641.25 179.36 642.96 ;
   RECT 0.00 642.96 179.36 644.67 ;
   RECT 0.00 644.67 179.36 646.38 ;
   RECT 0.00 646.38 179.36 648.09 ;
   RECT 0.00 648.09 179.36 649.80 ;
   RECT 0.00 649.80 179.36 651.51 ;
   RECT 0.00 651.51 179.36 653.22 ;
   RECT 0.00 653.22 179.36 654.93 ;
   RECT 0.00 654.93 179.36 656.64 ;
   RECT 0.00 656.64 179.36 658.35 ;
   RECT 0.00 658.35 179.36 660.06 ;
   RECT 0.00 660.06 179.36 661.77 ;
   RECT 0.00 661.77 179.36 663.48 ;
   RECT 0.00 663.48 179.36 665.19 ;
   RECT 0.00 665.19 179.36 666.90 ;
   RECT 0.00 666.90 179.36 668.61 ;
   RECT 0.00 668.61 179.36 670.32 ;
   RECT 0.00 670.32 179.36 672.03 ;
   RECT 0.00 672.03 179.36 673.74 ;
   RECT 0.00 673.74 179.36 675.45 ;
   RECT 0.00 675.45 179.36 677.16 ;
   RECT 0.00 677.16 179.36 678.87 ;
   RECT 0.00 678.87 179.36 680.58 ;
   RECT 0.00 680.58 179.36 682.29 ;
   RECT 0.00 682.29 179.36 684.00 ;
   RECT 0.00 684.00 179.36 685.71 ;
   RECT 0.00 685.71 179.36 687.42 ;
   RECT 0.00 687.42 179.36 689.13 ;
   RECT 0.00 689.13 179.36 690.84 ;
   RECT 0.00 690.84 179.36 692.55 ;
   RECT 0.00 692.55 179.36 694.26 ;
   RECT 0.00 694.26 179.36 695.97 ;
   RECT 0.00 695.97 179.36 697.68 ;
   RECT 0.00 697.68 179.36 699.39 ;
   RECT 0.00 699.39 179.36 701.10 ;
   RECT 0.00 701.10 179.36 702.81 ;
   RECT 0.00 702.81 179.36 704.52 ;
   RECT 0.00 704.52 179.36 706.23 ;
   RECT 0.00 706.23 179.36 707.94 ;
   RECT 0.00 707.94 179.36 709.65 ;
   RECT 0.00 709.65 179.36 711.36 ;
   RECT 0.00 711.36 179.36 713.07 ;
   RECT 0.00 713.07 179.36 714.78 ;
   RECT 0.00 714.78 179.36 716.49 ;
   RECT 0.00 716.49 179.36 718.20 ;
   RECT 0.00 718.20 179.36 719.91 ;
   RECT 0.00 719.91 179.36 721.62 ;
   RECT 0.00 721.62 179.36 723.33 ;
   RECT 0.00 723.33 179.36 725.04 ;
   RECT 0.00 725.04 179.36 726.75 ;
   RECT 0.00 726.75 179.36 728.46 ;
   RECT 0.00 728.46 179.36 730.17 ;
   RECT 0.00 730.17 179.36 731.88 ;
   RECT 0.00 731.88 179.36 733.59 ;
   RECT 0.00 733.59 179.36 735.30 ;
   RECT 0.00 735.30 179.36 737.01 ;
   RECT 0.00 737.01 179.36 738.72 ;
   RECT 0.00 738.72 179.36 740.43 ;
   RECT 0.00 740.43 179.36 742.14 ;
   RECT 0.00 742.14 179.36 743.85 ;
   RECT 0.00 743.85 179.36 745.56 ;
   RECT 0.00 745.56 179.36 747.27 ;
   RECT 0.00 747.27 179.36 748.98 ;
   RECT 0.00 748.98 179.36 750.69 ;
   RECT 0.00 750.69 179.36 752.40 ;
   RECT 0.00 752.40 179.36 754.11 ;
   RECT 0.00 754.11 179.36 755.82 ;
   RECT 0.00 755.82 179.36 757.53 ;
   RECT 0.00 757.53 179.36 759.24 ;
   RECT 0.00 759.24 179.36 760.95 ;
   RECT 0.00 760.95 179.36 762.66 ;
   RECT 0.00 762.66 179.36 764.37 ;
   RECT 0.00 764.37 179.36 766.08 ;
   RECT 0.00 766.08 179.36 767.79 ;
   RECT 0.00 767.79 179.36 769.50 ;
   RECT 0.00 769.50 179.36 771.21 ;
   RECT 0.00 771.21 179.36 772.92 ;
   RECT 0.00 772.92 179.36 774.63 ;
   RECT 0.00 774.63 179.36 776.34 ;
   RECT 0.00 776.34 179.36 778.05 ;
   RECT 0.00 778.05 179.36 779.76 ;
   RECT 0.00 779.76 179.36 781.47 ;
   RECT 0.00 781.47 179.36 783.18 ;
   RECT 0.00 783.18 179.36 784.89 ;
   RECT 0.00 784.89 179.36 786.60 ;
   RECT 0.00 786.60 179.36 788.31 ;
   RECT 0.00 788.31 179.36 790.02 ;
   RECT 0.00 790.02 179.36 791.73 ;
   RECT 0.00 791.73 179.36 793.44 ;
   RECT 0.00 793.44 179.36 795.15 ;
   RECT 0.00 795.15 179.36 796.86 ;
   RECT 0.00 796.86 179.36 798.57 ;
   RECT 0.00 798.57 179.36 800.28 ;
   RECT 0.00 800.28 179.36 801.99 ;
   RECT 0.00 801.99 179.36 803.70 ;
   RECT 0.00 803.70 179.36 805.41 ;
   RECT 0.00 805.41 179.36 807.12 ;
   RECT 0.00 807.12 179.36 808.83 ;
   RECT 0.00 808.83 179.36 810.54 ;
   RECT 0.00 810.54 179.36 812.25 ;
   RECT 0.00 812.25 179.36 813.96 ;
   RECT 0.00 813.96 179.36 815.67 ;
   RECT 0.00 815.67 179.36 817.38 ;
   RECT 0.00 817.38 179.36 819.09 ;
   RECT 0.00 819.09 179.36 820.80 ;
   RECT 0.00 820.80 179.36 822.51 ;
   RECT 0.00 822.51 179.36 824.22 ;
   RECT 0.00 824.22 179.36 825.93 ;
   RECT 0.00 825.93 179.36 827.64 ;
   RECT 0.00 827.64 179.36 829.35 ;
   RECT 0.00 829.35 179.36 831.06 ;
   RECT 0.00 831.06 179.36 832.77 ;
   RECT 0.00 832.77 179.36 834.48 ;
   RECT 0.00 834.48 179.36 836.19 ;
   RECT 0.00 836.19 179.36 837.90 ;
   RECT 0.00 837.90 179.36 839.61 ;
   RECT 0.00 839.61 179.36 841.32 ;
  LAYER via2 ;
   RECT 0.00 0.00 179.36 1.71 ;
   RECT 0.00 1.71 179.36 3.42 ;
   RECT 0.00 3.42 179.36 5.13 ;
   RECT 0.00 5.13 179.36 6.84 ;
   RECT 0.00 6.84 179.36 8.55 ;
   RECT 0.00 8.55 179.36 10.26 ;
   RECT 0.00 10.26 179.36 11.97 ;
   RECT 0.00 11.97 179.36 13.68 ;
   RECT 0.00 13.68 179.36 15.39 ;
   RECT 0.00 15.39 179.36 17.10 ;
   RECT 0.00 17.10 179.36 18.81 ;
   RECT 0.00 18.81 179.36 20.52 ;
   RECT 0.00 20.52 179.36 22.23 ;
   RECT 0.00 22.23 179.36 23.94 ;
   RECT 0.00 23.94 179.36 25.65 ;
   RECT 0.00 25.65 179.36 27.36 ;
   RECT 0.00 27.36 179.36 29.07 ;
   RECT 0.00 29.07 179.36 30.78 ;
   RECT 0.00 30.78 179.36 32.49 ;
   RECT 0.00 32.49 179.36 34.20 ;
   RECT 0.00 34.20 179.36 35.91 ;
   RECT 0.00 35.91 179.36 37.62 ;
   RECT 0.00 37.62 179.36 39.33 ;
   RECT 0.00 39.33 179.36 41.04 ;
   RECT 0.00 41.04 179.36 42.75 ;
   RECT 0.00 42.75 179.36 44.46 ;
   RECT 0.00 44.46 179.36 46.17 ;
   RECT 0.00 46.17 179.36 47.88 ;
   RECT 0.00 47.88 179.36 49.59 ;
   RECT 0.00 49.59 179.36 51.30 ;
   RECT 0.00 51.30 179.36 53.01 ;
   RECT 0.00 53.01 179.36 54.72 ;
   RECT 0.00 54.72 179.36 56.43 ;
   RECT 0.00 56.43 179.36 58.14 ;
   RECT 0.00 58.14 179.36 59.85 ;
   RECT 0.00 59.85 179.36 61.56 ;
   RECT 0.00 61.56 179.36 63.27 ;
   RECT 0.00 63.27 179.36 64.98 ;
   RECT 0.00 64.98 179.36 66.69 ;
   RECT 0.00 66.69 179.36 68.40 ;
   RECT 0.00 68.40 179.36 70.11 ;
   RECT 0.00 70.11 179.36 71.82 ;
   RECT 0.00 71.82 179.36 73.53 ;
   RECT 0.00 73.53 179.36 75.24 ;
   RECT 0.00 75.24 179.36 76.95 ;
   RECT 0.00 76.95 179.36 78.66 ;
   RECT 0.00 78.66 179.36 80.37 ;
   RECT 0.00 80.37 179.36 82.08 ;
   RECT 0.00 82.08 179.36 83.79 ;
   RECT 0.00 83.79 179.36 85.50 ;
   RECT 0.00 85.50 179.36 87.21 ;
   RECT 0.00 87.21 179.36 88.92 ;
   RECT 0.00 88.92 179.36 90.63 ;
   RECT 0.00 90.63 179.36 92.34 ;
   RECT 0.00 92.34 179.36 94.05 ;
   RECT 0.00 94.05 179.36 95.76 ;
   RECT 0.00 95.76 179.36 97.47 ;
   RECT 0.00 97.47 179.36 99.18 ;
   RECT 0.00 99.18 179.36 100.89 ;
   RECT 0.00 100.89 179.36 102.60 ;
   RECT 0.00 102.60 179.36 104.31 ;
   RECT 0.00 104.31 179.36 106.02 ;
   RECT 0.00 106.02 179.36 107.73 ;
   RECT 0.00 107.73 179.36 109.44 ;
   RECT 0.00 109.44 179.36 111.15 ;
   RECT 0.00 111.15 179.36 112.86 ;
   RECT 0.00 112.86 179.36 114.57 ;
   RECT 0.00 114.57 179.36 116.28 ;
   RECT 0.00 116.28 179.36 117.99 ;
   RECT 0.00 117.99 179.36 119.70 ;
   RECT 0.00 119.70 179.36 121.41 ;
   RECT 0.00 121.41 179.36 123.12 ;
   RECT 0.00 123.12 179.36 124.83 ;
   RECT 0.00 124.83 179.36 126.54 ;
   RECT 0.00 126.54 179.36 128.25 ;
   RECT 0.00 128.25 179.36 129.96 ;
   RECT 0.00 129.96 179.36 131.67 ;
   RECT 0.00 131.67 179.36 133.38 ;
   RECT 0.00 133.38 179.36 135.09 ;
   RECT 0.00 135.09 179.36 136.80 ;
   RECT 0.00 136.80 179.36 138.51 ;
   RECT 0.00 138.51 179.36 140.22 ;
   RECT 0.00 140.22 179.36 141.93 ;
   RECT 0.00 141.93 179.36 143.64 ;
   RECT 0.00 143.64 179.36 145.35 ;
   RECT 0.00 145.35 179.36 147.06 ;
   RECT 0.00 147.06 179.36 148.77 ;
   RECT 0.00 148.77 179.36 150.48 ;
   RECT 0.00 150.48 179.36 152.19 ;
   RECT 0.00 152.19 179.36 153.90 ;
   RECT 0.00 153.90 179.36 155.61 ;
   RECT 0.00 155.61 179.36 157.32 ;
   RECT 0.00 157.32 179.36 159.03 ;
   RECT 0.00 159.03 179.36 160.74 ;
   RECT 0.00 160.74 179.36 162.45 ;
   RECT 0.00 162.45 179.36 164.16 ;
   RECT 0.00 164.16 179.36 165.87 ;
   RECT 0.00 165.87 179.36 167.58 ;
   RECT 0.00 167.58 179.36 169.29 ;
   RECT 0.00 169.29 179.36 171.00 ;
   RECT 0.00 171.00 179.36 172.71 ;
   RECT 0.00 172.71 179.36 174.42 ;
   RECT 0.00 174.42 179.36 176.13 ;
   RECT 0.00 176.13 179.36 177.84 ;
   RECT 0.00 177.84 179.36 179.55 ;
   RECT 0.00 179.55 179.36 181.26 ;
   RECT 0.00 181.26 179.36 182.97 ;
   RECT 0.00 182.97 179.36 184.68 ;
   RECT 0.00 184.68 179.36 186.39 ;
   RECT 0.00 186.39 179.36 188.10 ;
   RECT 0.00 188.10 179.36 189.81 ;
   RECT 0.00 189.81 179.36 191.52 ;
   RECT 0.00 191.52 179.36 193.23 ;
   RECT 0.00 193.23 179.36 194.94 ;
   RECT 0.00 194.94 179.36 196.65 ;
   RECT 0.00 196.65 179.36 198.36 ;
   RECT 0.00 198.36 179.36 200.07 ;
   RECT 0.00 200.07 179.36 201.78 ;
   RECT 0.00 201.78 179.36 203.49 ;
   RECT 0.00 203.49 179.36 205.20 ;
   RECT 0.00 205.20 179.36 206.91 ;
   RECT 0.00 206.91 179.36 208.62 ;
   RECT 0.00 208.62 179.36 210.33 ;
   RECT 0.00 210.33 179.36 212.04 ;
   RECT 0.00 212.04 179.36 213.75 ;
   RECT 0.00 213.75 179.36 215.46 ;
   RECT 0.00 215.46 179.36 217.17 ;
   RECT 0.00 217.17 179.36 218.88 ;
   RECT 0.00 218.88 179.36 220.59 ;
   RECT 0.00 220.59 179.36 222.30 ;
   RECT 0.00 222.30 179.36 224.01 ;
   RECT 0.00 224.01 179.36 225.72 ;
   RECT 0.00 225.72 179.36 227.43 ;
   RECT 0.00 227.43 179.36 229.14 ;
   RECT 0.00 229.14 179.36 230.85 ;
   RECT 0.00 230.85 179.36 232.56 ;
   RECT 0.00 232.56 179.36 234.27 ;
   RECT 0.00 234.27 179.36 235.98 ;
   RECT 0.00 235.98 179.36 237.69 ;
   RECT 0.00 237.69 179.36 239.40 ;
   RECT 0.00 239.40 179.36 241.11 ;
   RECT 0.00 241.11 179.36 242.82 ;
   RECT 0.00 242.82 179.36 244.53 ;
   RECT 0.00 244.53 179.36 246.24 ;
   RECT 0.00 246.24 179.36 247.95 ;
   RECT 0.00 247.95 179.36 249.66 ;
   RECT 0.00 249.66 179.36 251.37 ;
   RECT 0.00 251.37 179.36 253.08 ;
   RECT 0.00 253.08 179.36 254.79 ;
   RECT 0.00 254.79 179.36 256.50 ;
   RECT 0.00 256.50 179.36 258.21 ;
   RECT 0.00 258.21 179.36 259.92 ;
   RECT 0.00 259.92 179.36 261.63 ;
   RECT 0.00 261.63 179.36 263.34 ;
   RECT 0.00 263.34 179.36 265.05 ;
   RECT 0.00 265.05 179.36 266.76 ;
   RECT 0.00 266.76 179.36 268.47 ;
   RECT 0.00 268.47 179.36 270.18 ;
   RECT 0.00 270.18 179.36 271.89 ;
   RECT 0.00 271.89 179.36 273.60 ;
   RECT 0.00 273.60 179.36 275.31 ;
   RECT 0.00 275.31 179.36 277.02 ;
   RECT 0.00 277.02 179.36 278.73 ;
   RECT 0.00 278.73 179.36 280.44 ;
   RECT 0.00 280.44 179.36 282.15 ;
   RECT 0.00 282.15 179.36 283.86 ;
   RECT 0.00 283.86 179.36 285.57 ;
   RECT 0.00 285.57 179.36 287.28 ;
   RECT 0.00 287.28 179.36 288.99 ;
   RECT 0.00 288.99 179.36 290.70 ;
   RECT 0.00 290.70 179.36 292.41 ;
   RECT 0.00 292.41 179.36 294.12 ;
   RECT 0.00 294.12 179.36 295.83 ;
   RECT 0.00 295.83 179.36 297.54 ;
   RECT 0.00 297.54 179.36 299.25 ;
   RECT 0.00 299.25 179.36 300.96 ;
   RECT 0.00 300.96 179.36 302.67 ;
   RECT 0.00 302.67 179.36 304.38 ;
   RECT 0.00 304.38 179.36 306.09 ;
   RECT 0.00 306.09 179.36 307.80 ;
   RECT 0.00 307.80 179.36 309.51 ;
   RECT 0.00 309.51 179.36 311.22 ;
   RECT 0.00 311.22 179.36 312.93 ;
   RECT 0.00 312.93 179.36 314.64 ;
   RECT 0.00 314.64 179.36 316.35 ;
   RECT 0.00 316.35 179.36 318.06 ;
   RECT 0.00 318.06 179.36 319.77 ;
   RECT 0.00 319.77 179.36 321.48 ;
   RECT 0.00 321.48 179.36 323.19 ;
   RECT 0.00 323.19 179.36 324.90 ;
   RECT 0.00 324.90 179.36 326.61 ;
   RECT 0.00 326.61 179.36 328.32 ;
   RECT 0.00 328.32 179.36 330.03 ;
   RECT 0.00 330.03 179.36 331.74 ;
   RECT 0.00 331.74 179.36 333.45 ;
   RECT 0.00 333.45 179.36 335.16 ;
   RECT 0.00 335.16 179.36 336.87 ;
   RECT 0.00 336.87 179.36 338.58 ;
   RECT 0.00 338.58 179.36 340.29 ;
   RECT 0.00 340.29 179.36 342.00 ;
   RECT 0.00 342.00 179.36 343.71 ;
   RECT 0.00 343.71 179.36 345.42 ;
   RECT 0.00 345.42 179.36 347.13 ;
   RECT 0.00 347.13 179.36 348.84 ;
   RECT 0.00 348.84 179.36 350.55 ;
   RECT 0.00 350.55 179.36 352.26 ;
   RECT 0.00 352.26 179.36 353.97 ;
   RECT 0.00 353.97 179.36 355.68 ;
   RECT 0.00 355.68 179.36 357.39 ;
   RECT 0.00 357.39 179.36 359.10 ;
   RECT 0.00 359.10 179.36 360.81 ;
   RECT 0.00 360.81 179.36 362.52 ;
   RECT 0.00 362.52 179.36 364.23 ;
   RECT 0.00 364.23 179.36 365.94 ;
   RECT 0.00 365.94 179.36 367.65 ;
   RECT 0.00 367.65 179.36 369.36 ;
   RECT 0.00 369.36 179.36 371.07 ;
   RECT 0.00 371.07 179.36 372.78 ;
   RECT 0.00 372.78 179.36 374.49 ;
   RECT 0.00 374.49 179.36 376.20 ;
   RECT 0.00 376.20 179.36 377.91 ;
   RECT 0.00 377.91 179.36 379.62 ;
   RECT 0.00 379.62 179.36 381.33 ;
   RECT 0.00 381.33 179.36 383.04 ;
   RECT 0.00 383.04 179.36 384.75 ;
   RECT 0.00 384.75 179.36 386.46 ;
   RECT 0.00 386.46 179.36 388.17 ;
   RECT 0.00 388.17 179.36 389.88 ;
   RECT 0.00 389.88 179.36 391.59 ;
   RECT 0.00 391.59 179.36 393.30 ;
   RECT 0.00 393.30 179.36 395.01 ;
   RECT 0.00 395.01 179.36 396.72 ;
   RECT 0.00 396.72 179.36 398.43 ;
   RECT 0.00 398.43 179.36 400.14 ;
   RECT 0.00 400.14 179.36 401.85 ;
   RECT 0.00 401.85 202.54 403.56 ;
   RECT 0.00 403.56 202.54 405.27 ;
   RECT 0.00 405.27 202.54 406.98 ;
   RECT 0.00 406.98 202.54 408.69 ;
   RECT 0.00 408.69 202.54 410.40 ;
   RECT 0.00 410.40 202.54 412.11 ;
   RECT 0.00 412.11 202.54 413.82 ;
   RECT 0.00 413.82 202.54 415.53 ;
   RECT 0.00 415.53 202.54 417.24 ;
   RECT 0.00 417.24 202.54 418.95 ;
   RECT 0.00 418.95 202.54 420.66 ;
   RECT 0.00 420.66 202.54 422.37 ;
   RECT 0.00 422.37 202.54 424.08 ;
   RECT 0.00 424.08 202.54 425.79 ;
   RECT 0.00 425.79 202.54 427.50 ;
   RECT 0.00 427.50 202.54 429.21 ;
   RECT 0.00 429.21 202.54 430.92 ;
   RECT 0.00 430.92 179.36 432.63 ;
   RECT 0.00 432.63 179.36 434.34 ;
   RECT 0.00 434.34 179.36 436.05 ;
   RECT 0.00 436.05 179.36 437.76 ;
   RECT 0.00 437.76 179.36 439.47 ;
   RECT 0.00 439.47 179.36 441.18 ;
   RECT 0.00 441.18 179.36 442.89 ;
   RECT 0.00 442.89 179.36 444.60 ;
   RECT 0.00 444.60 179.36 446.31 ;
   RECT 0.00 446.31 179.36 448.02 ;
   RECT 0.00 448.02 179.36 449.73 ;
   RECT 0.00 449.73 179.36 451.44 ;
   RECT 0.00 451.44 179.36 453.15 ;
   RECT 0.00 453.15 179.36 454.86 ;
   RECT 0.00 454.86 179.36 456.57 ;
   RECT 0.00 456.57 179.36 458.28 ;
   RECT 0.00 458.28 179.36 459.99 ;
   RECT 0.00 459.99 179.36 461.70 ;
   RECT 0.00 461.70 179.36 463.41 ;
   RECT 0.00 463.41 179.36 465.12 ;
   RECT 0.00 465.12 179.36 466.83 ;
   RECT 0.00 466.83 179.36 468.54 ;
   RECT 0.00 468.54 179.36 470.25 ;
   RECT 0.00 470.25 179.36 471.96 ;
   RECT 0.00 471.96 179.36 473.67 ;
   RECT 0.00 473.67 179.36 475.38 ;
   RECT 0.00 475.38 179.36 477.09 ;
   RECT 0.00 477.09 179.36 478.80 ;
   RECT 0.00 478.80 179.36 480.51 ;
   RECT 0.00 480.51 179.36 482.22 ;
   RECT 0.00 482.22 179.36 483.93 ;
   RECT 0.00 483.93 179.36 485.64 ;
   RECT 0.00 485.64 179.36 487.35 ;
   RECT 0.00 487.35 179.36 489.06 ;
   RECT 0.00 489.06 179.36 490.77 ;
   RECT 0.00 490.77 179.36 492.48 ;
   RECT 0.00 492.48 179.36 494.19 ;
   RECT 0.00 494.19 179.36 495.90 ;
   RECT 0.00 495.90 179.36 497.61 ;
   RECT 0.00 497.61 179.36 499.32 ;
   RECT 0.00 499.32 179.36 501.03 ;
   RECT 0.00 501.03 179.36 502.74 ;
   RECT 0.00 502.74 179.36 504.45 ;
   RECT 0.00 504.45 179.36 506.16 ;
   RECT 0.00 506.16 179.36 507.87 ;
   RECT 0.00 507.87 179.36 509.58 ;
   RECT 0.00 509.58 179.36 511.29 ;
   RECT 0.00 511.29 179.36 513.00 ;
   RECT 0.00 513.00 179.36 514.71 ;
   RECT 0.00 514.71 179.36 516.42 ;
   RECT 0.00 516.42 179.36 518.13 ;
   RECT 0.00 518.13 179.36 519.84 ;
   RECT 0.00 519.84 179.36 521.55 ;
   RECT 0.00 521.55 179.36 523.26 ;
   RECT 0.00 523.26 179.36 524.97 ;
   RECT 0.00 524.97 179.36 526.68 ;
   RECT 0.00 526.68 179.36 528.39 ;
   RECT 0.00 528.39 179.36 530.10 ;
   RECT 0.00 530.10 179.36 531.81 ;
   RECT 0.00 531.81 179.36 533.52 ;
   RECT 0.00 533.52 179.36 535.23 ;
   RECT 0.00 535.23 179.36 536.94 ;
   RECT 0.00 536.94 179.36 538.65 ;
   RECT 0.00 538.65 179.36 540.36 ;
   RECT 0.00 540.36 179.36 542.07 ;
   RECT 0.00 542.07 179.36 543.78 ;
   RECT 0.00 543.78 179.36 545.49 ;
   RECT 0.00 545.49 179.36 547.20 ;
   RECT 0.00 547.20 179.36 548.91 ;
   RECT 0.00 548.91 179.36 550.62 ;
   RECT 0.00 550.62 179.36 552.33 ;
   RECT 0.00 552.33 179.36 554.04 ;
   RECT 0.00 554.04 179.36 555.75 ;
   RECT 0.00 555.75 179.36 557.46 ;
   RECT 0.00 557.46 179.36 559.17 ;
   RECT 0.00 559.17 179.36 560.88 ;
   RECT 0.00 560.88 179.36 562.59 ;
   RECT 0.00 562.59 179.36 564.30 ;
   RECT 0.00 564.30 179.36 566.01 ;
   RECT 0.00 566.01 179.36 567.72 ;
   RECT 0.00 567.72 179.36 569.43 ;
   RECT 0.00 569.43 179.36 571.14 ;
   RECT 0.00 571.14 179.36 572.85 ;
   RECT 0.00 572.85 179.36 574.56 ;
   RECT 0.00 574.56 179.36 576.27 ;
   RECT 0.00 576.27 179.36 577.98 ;
   RECT 0.00 577.98 179.36 579.69 ;
   RECT 0.00 579.69 179.36 581.40 ;
   RECT 0.00 581.40 179.36 583.11 ;
   RECT 0.00 583.11 179.36 584.82 ;
   RECT 0.00 584.82 179.36 586.53 ;
   RECT 0.00 586.53 179.36 588.24 ;
   RECT 0.00 588.24 179.36 589.95 ;
   RECT 0.00 589.95 179.36 591.66 ;
   RECT 0.00 591.66 179.36 593.37 ;
   RECT 0.00 593.37 179.36 595.08 ;
   RECT 0.00 595.08 179.36 596.79 ;
   RECT 0.00 596.79 179.36 598.50 ;
   RECT 0.00 598.50 179.36 600.21 ;
   RECT 0.00 600.21 179.36 601.92 ;
   RECT 0.00 601.92 179.36 603.63 ;
   RECT 0.00 603.63 179.36 605.34 ;
   RECT 0.00 605.34 179.36 607.05 ;
   RECT 0.00 607.05 179.36 608.76 ;
   RECT 0.00 608.76 179.36 610.47 ;
   RECT 0.00 610.47 179.36 612.18 ;
   RECT 0.00 612.18 179.36 613.89 ;
   RECT 0.00 613.89 179.36 615.60 ;
   RECT 0.00 615.60 179.36 617.31 ;
   RECT 0.00 617.31 179.36 619.02 ;
   RECT 0.00 619.02 179.36 620.73 ;
   RECT 0.00 620.73 179.36 622.44 ;
   RECT 0.00 622.44 179.36 624.15 ;
   RECT 0.00 624.15 179.36 625.86 ;
   RECT 0.00 625.86 179.36 627.57 ;
   RECT 0.00 627.57 179.36 629.28 ;
   RECT 0.00 629.28 179.36 630.99 ;
   RECT 0.00 630.99 179.36 632.70 ;
   RECT 0.00 632.70 179.36 634.41 ;
   RECT 0.00 634.41 179.36 636.12 ;
   RECT 0.00 636.12 179.36 637.83 ;
   RECT 0.00 637.83 179.36 639.54 ;
   RECT 0.00 639.54 179.36 641.25 ;
   RECT 0.00 641.25 179.36 642.96 ;
   RECT 0.00 642.96 179.36 644.67 ;
   RECT 0.00 644.67 179.36 646.38 ;
   RECT 0.00 646.38 179.36 648.09 ;
   RECT 0.00 648.09 179.36 649.80 ;
   RECT 0.00 649.80 179.36 651.51 ;
   RECT 0.00 651.51 179.36 653.22 ;
   RECT 0.00 653.22 179.36 654.93 ;
   RECT 0.00 654.93 179.36 656.64 ;
   RECT 0.00 656.64 179.36 658.35 ;
   RECT 0.00 658.35 179.36 660.06 ;
   RECT 0.00 660.06 179.36 661.77 ;
   RECT 0.00 661.77 179.36 663.48 ;
   RECT 0.00 663.48 179.36 665.19 ;
   RECT 0.00 665.19 179.36 666.90 ;
   RECT 0.00 666.90 179.36 668.61 ;
   RECT 0.00 668.61 179.36 670.32 ;
   RECT 0.00 670.32 179.36 672.03 ;
   RECT 0.00 672.03 179.36 673.74 ;
   RECT 0.00 673.74 179.36 675.45 ;
   RECT 0.00 675.45 179.36 677.16 ;
   RECT 0.00 677.16 179.36 678.87 ;
   RECT 0.00 678.87 179.36 680.58 ;
   RECT 0.00 680.58 179.36 682.29 ;
   RECT 0.00 682.29 179.36 684.00 ;
   RECT 0.00 684.00 179.36 685.71 ;
   RECT 0.00 685.71 179.36 687.42 ;
   RECT 0.00 687.42 179.36 689.13 ;
   RECT 0.00 689.13 179.36 690.84 ;
   RECT 0.00 690.84 179.36 692.55 ;
   RECT 0.00 692.55 179.36 694.26 ;
   RECT 0.00 694.26 179.36 695.97 ;
   RECT 0.00 695.97 179.36 697.68 ;
   RECT 0.00 697.68 179.36 699.39 ;
   RECT 0.00 699.39 179.36 701.10 ;
   RECT 0.00 701.10 179.36 702.81 ;
   RECT 0.00 702.81 179.36 704.52 ;
   RECT 0.00 704.52 179.36 706.23 ;
   RECT 0.00 706.23 179.36 707.94 ;
   RECT 0.00 707.94 179.36 709.65 ;
   RECT 0.00 709.65 179.36 711.36 ;
   RECT 0.00 711.36 179.36 713.07 ;
   RECT 0.00 713.07 179.36 714.78 ;
   RECT 0.00 714.78 179.36 716.49 ;
   RECT 0.00 716.49 179.36 718.20 ;
   RECT 0.00 718.20 179.36 719.91 ;
   RECT 0.00 719.91 179.36 721.62 ;
   RECT 0.00 721.62 179.36 723.33 ;
   RECT 0.00 723.33 179.36 725.04 ;
   RECT 0.00 725.04 179.36 726.75 ;
   RECT 0.00 726.75 179.36 728.46 ;
   RECT 0.00 728.46 179.36 730.17 ;
   RECT 0.00 730.17 179.36 731.88 ;
   RECT 0.00 731.88 179.36 733.59 ;
   RECT 0.00 733.59 179.36 735.30 ;
   RECT 0.00 735.30 179.36 737.01 ;
   RECT 0.00 737.01 179.36 738.72 ;
   RECT 0.00 738.72 179.36 740.43 ;
   RECT 0.00 740.43 179.36 742.14 ;
   RECT 0.00 742.14 179.36 743.85 ;
   RECT 0.00 743.85 179.36 745.56 ;
   RECT 0.00 745.56 179.36 747.27 ;
   RECT 0.00 747.27 179.36 748.98 ;
   RECT 0.00 748.98 179.36 750.69 ;
   RECT 0.00 750.69 179.36 752.40 ;
   RECT 0.00 752.40 179.36 754.11 ;
   RECT 0.00 754.11 179.36 755.82 ;
   RECT 0.00 755.82 179.36 757.53 ;
   RECT 0.00 757.53 179.36 759.24 ;
   RECT 0.00 759.24 179.36 760.95 ;
   RECT 0.00 760.95 179.36 762.66 ;
   RECT 0.00 762.66 179.36 764.37 ;
   RECT 0.00 764.37 179.36 766.08 ;
   RECT 0.00 766.08 179.36 767.79 ;
   RECT 0.00 767.79 179.36 769.50 ;
   RECT 0.00 769.50 179.36 771.21 ;
   RECT 0.00 771.21 179.36 772.92 ;
   RECT 0.00 772.92 179.36 774.63 ;
   RECT 0.00 774.63 179.36 776.34 ;
   RECT 0.00 776.34 179.36 778.05 ;
   RECT 0.00 778.05 179.36 779.76 ;
   RECT 0.00 779.76 179.36 781.47 ;
   RECT 0.00 781.47 179.36 783.18 ;
   RECT 0.00 783.18 179.36 784.89 ;
   RECT 0.00 784.89 179.36 786.60 ;
   RECT 0.00 786.60 179.36 788.31 ;
   RECT 0.00 788.31 179.36 790.02 ;
   RECT 0.00 790.02 179.36 791.73 ;
   RECT 0.00 791.73 179.36 793.44 ;
   RECT 0.00 793.44 179.36 795.15 ;
   RECT 0.00 795.15 179.36 796.86 ;
   RECT 0.00 796.86 179.36 798.57 ;
   RECT 0.00 798.57 179.36 800.28 ;
   RECT 0.00 800.28 179.36 801.99 ;
   RECT 0.00 801.99 179.36 803.70 ;
   RECT 0.00 803.70 179.36 805.41 ;
   RECT 0.00 805.41 179.36 807.12 ;
   RECT 0.00 807.12 179.36 808.83 ;
   RECT 0.00 808.83 179.36 810.54 ;
   RECT 0.00 810.54 179.36 812.25 ;
   RECT 0.00 812.25 179.36 813.96 ;
   RECT 0.00 813.96 179.36 815.67 ;
   RECT 0.00 815.67 179.36 817.38 ;
   RECT 0.00 817.38 179.36 819.09 ;
   RECT 0.00 819.09 179.36 820.80 ;
   RECT 0.00 820.80 179.36 822.51 ;
   RECT 0.00 822.51 179.36 824.22 ;
   RECT 0.00 824.22 179.36 825.93 ;
   RECT 0.00 825.93 179.36 827.64 ;
   RECT 0.00 827.64 179.36 829.35 ;
   RECT 0.00 829.35 179.36 831.06 ;
   RECT 0.00 831.06 179.36 832.77 ;
   RECT 0.00 832.77 179.36 834.48 ;
   RECT 0.00 834.48 179.36 836.19 ;
   RECT 0.00 836.19 179.36 837.90 ;
   RECT 0.00 837.90 179.36 839.61 ;
   RECT 0.00 839.61 179.36 841.32 ;
  LAYER metal3 ;
   RECT 0.00 0.00 179.36 1.71 ;
   RECT 0.00 1.71 179.36 3.42 ;
   RECT 0.00 3.42 179.36 5.13 ;
   RECT 0.00 5.13 179.36 6.84 ;
   RECT 0.00 6.84 179.36 8.55 ;
   RECT 0.00 8.55 179.36 10.26 ;
   RECT 0.00 10.26 179.36 11.97 ;
   RECT 0.00 11.97 179.36 13.68 ;
   RECT 0.00 13.68 179.36 15.39 ;
   RECT 0.00 15.39 179.36 17.10 ;
   RECT 0.00 17.10 179.36 18.81 ;
   RECT 0.00 18.81 179.36 20.52 ;
   RECT 0.00 20.52 179.36 22.23 ;
   RECT 0.00 22.23 179.36 23.94 ;
   RECT 0.00 23.94 179.36 25.65 ;
   RECT 0.00 25.65 179.36 27.36 ;
   RECT 0.00 27.36 179.36 29.07 ;
   RECT 0.00 29.07 179.36 30.78 ;
   RECT 0.00 30.78 179.36 32.49 ;
   RECT 0.00 32.49 179.36 34.20 ;
   RECT 0.00 34.20 179.36 35.91 ;
   RECT 0.00 35.91 179.36 37.62 ;
   RECT 0.00 37.62 179.36 39.33 ;
   RECT 0.00 39.33 179.36 41.04 ;
   RECT 0.00 41.04 179.36 42.75 ;
   RECT 0.00 42.75 179.36 44.46 ;
   RECT 0.00 44.46 179.36 46.17 ;
   RECT 0.00 46.17 179.36 47.88 ;
   RECT 0.00 47.88 179.36 49.59 ;
   RECT 0.00 49.59 179.36 51.30 ;
   RECT 0.00 51.30 179.36 53.01 ;
   RECT 0.00 53.01 179.36 54.72 ;
   RECT 0.00 54.72 179.36 56.43 ;
   RECT 0.00 56.43 179.36 58.14 ;
   RECT 0.00 58.14 179.36 59.85 ;
   RECT 0.00 59.85 179.36 61.56 ;
   RECT 0.00 61.56 179.36 63.27 ;
   RECT 0.00 63.27 179.36 64.98 ;
   RECT 0.00 64.98 179.36 66.69 ;
   RECT 0.00 66.69 179.36 68.40 ;
   RECT 0.00 68.40 179.36 70.11 ;
   RECT 0.00 70.11 179.36 71.82 ;
   RECT 0.00 71.82 179.36 73.53 ;
   RECT 0.00 73.53 179.36 75.24 ;
   RECT 0.00 75.24 179.36 76.95 ;
   RECT 0.00 76.95 179.36 78.66 ;
   RECT 0.00 78.66 179.36 80.37 ;
   RECT 0.00 80.37 179.36 82.08 ;
   RECT 0.00 82.08 179.36 83.79 ;
   RECT 0.00 83.79 179.36 85.50 ;
   RECT 0.00 85.50 179.36 87.21 ;
   RECT 0.00 87.21 179.36 88.92 ;
   RECT 0.00 88.92 179.36 90.63 ;
   RECT 0.00 90.63 179.36 92.34 ;
   RECT 0.00 92.34 179.36 94.05 ;
   RECT 0.00 94.05 179.36 95.76 ;
   RECT 0.00 95.76 179.36 97.47 ;
   RECT 0.00 97.47 179.36 99.18 ;
   RECT 0.00 99.18 179.36 100.89 ;
   RECT 0.00 100.89 179.36 102.60 ;
   RECT 0.00 102.60 179.36 104.31 ;
   RECT 0.00 104.31 179.36 106.02 ;
   RECT 0.00 106.02 179.36 107.73 ;
   RECT 0.00 107.73 179.36 109.44 ;
   RECT 0.00 109.44 179.36 111.15 ;
   RECT 0.00 111.15 179.36 112.86 ;
   RECT 0.00 112.86 179.36 114.57 ;
   RECT 0.00 114.57 179.36 116.28 ;
   RECT 0.00 116.28 179.36 117.99 ;
   RECT 0.00 117.99 179.36 119.70 ;
   RECT 0.00 119.70 179.36 121.41 ;
   RECT 0.00 121.41 179.36 123.12 ;
   RECT 0.00 123.12 179.36 124.83 ;
   RECT 0.00 124.83 179.36 126.54 ;
   RECT 0.00 126.54 179.36 128.25 ;
   RECT 0.00 128.25 179.36 129.96 ;
   RECT 0.00 129.96 179.36 131.67 ;
   RECT 0.00 131.67 179.36 133.38 ;
   RECT 0.00 133.38 179.36 135.09 ;
   RECT 0.00 135.09 179.36 136.80 ;
   RECT 0.00 136.80 179.36 138.51 ;
   RECT 0.00 138.51 179.36 140.22 ;
   RECT 0.00 140.22 179.36 141.93 ;
   RECT 0.00 141.93 179.36 143.64 ;
   RECT 0.00 143.64 179.36 145.35 ;
   RECT 0.00 145.35 179.36 147.06 ;
   RECT 0.00 147.06 179.36 148.77 ;
   RECT 0.00 148.77 179.36 150.48 ;
   RECT 0.00 150.48 179.36 152.19 ;
   RECT 0.00 152.19 179.36 153.90 ;
   RECT 0.00 153.90 179.36 155.61 ;
   RECT 0.00 155.61 179.36 157.32 ;
   RECT 0.00 157.32 179.36 159.03 ;
   RECT 0.00 159.03 179.36 160.74 ;
   RECT 0.00 160.74 179.36 162.45 ;
   RECT 0.00 162.45 179.36 164.16 ;
   RECT 0.00 164.16 179.36 165.87 ;
   RECT 0.00 165.87 179.36 167.58 ;
   RECT 0.00 167.58 179.36 169.29 ;
   RECT 0.00 169.29 179.36 171.00 ;
   RECT 0.00 171.00 179.36 172.71 ;
   RECT 0.00 172.71 179.36 174.42 ;
   RECT 0.00 174.42 179.36 176.13 ;
   RECT 0.00 176.13 179.36 177.84 ;
   RECT 0.00 177.84 179.36 179.55 ;
   RECT 0.00 179.55 179.36 181.26 ;
   RECT 0.00 181.26 179.36 182.97 ;
   RECT 0.00 182.97 179.36 184.68 ;
   RECT 0.00 184.68 179.36 186.39 ;
   RECT 0.00 186.39 179.36 188.10 ;
   RECT 0.00 188.10 179.36 189.81 ;
   RECT 0.00 189.81 179.36 191.52 ;
   RECT 0.00 191.52 179.36 193.23 ;
   RECT 0.00 193.23 179.36 194.94 ;
   RECT 0.00 194.94 179.36 196.65 ;
   RECT 0.00 196.65 179.36 198.36 ;
   RECT 0.00 198.36 179.36 200.07 ;
   RECT 0.00 200.07 179.36 201.78 ;
   RECT 0.00 201.78 179.36 203.49 ;
   RECT 0.00 203.49 179.36 205.20 ;
   RECT 0.00 205.20 179.36 206.91 ;
   RECT 0.00 206.91 179.36 208.62 ;
   RECT 0.00 208.62 179.36 210.33 ;
   RECT 0.00 210.33 179.36 212.04 ;
   RECT 0.00 212.04 179.36 213.75 ;
   RECT 0.00 213.75 179.36 215.46 ;
   RECT 0.00 215.46 179.36 217.17 ;
   RECT 0.00 217.17 179.36 218.88 ;
   RECT 0.00 218.88 179.36 220.59 ;
   RECT 0.00 220.59 179.36 222.30 ;
   RECT 0.00 222.30 179.36 224.01 ;
   RECT 0.00 224.01 179.36 225.72 ;
   RECT 0.00 225.72 179.36 227.43 ;
   RECT 0.00 227.43 179.36 229.14 ;
   RECT 0.00 229.14 179.36 230.85 ;
   RECT 0.00 230.85 179.36 232.56 ;
   RECT 0.00 232.56 179.36 234.27 ;
   RECT 0.00 234.27 179.36 235.98 ;
   RECT 0.00 235.98 179.36 237.69 ;
   RECT 0.00 237.69 179.36 239.40 ;
   RECT 0.00 239.40 179.36 241.11 ;
   RECT 0.00 241.11 179.36 242.82 ;
   RECT 0.00 242.82 179.36 244.53 ;
   RECT 0.00 244.53 179.36 246.24 ;
   RECT 0.00 246.24 179.36 247.95 ;
   RECT 0.00 247.95 179.36 249.66 ;
   RECT 0.00 249.66 179.36 251.37 ;
   RECT 0.00 251.37 179.36 253.08 ;
   RECT 0.00 253.08 179.36 254.79 ;
   RECT 0.00 254.79 179.36 256.50 ;
   RECT 0.00 256.50 179.36 258.21 ;
   RECT 0.00 258.21 179.36 259.92 ;
   RECT 0.00 259.92 179.36 261.63 ;
   RECT 0.00 261.63 179.36 263.34 ;
   RECT 0.00 263.34 179.36 265.05 ;
   RECT 0.00 265.05 179.36 266.76 ;
   RECT 0.00 266.76 179.36 268.47 ;
   RECT 0.00 268.47 179.36 270.18 ;
   RECT 0.00 270.18 179.36 271.89 ;
   RECT 0.00 271.89 179.36 273.60 ;
   RECT 0.00 273.60 179.36 275.31 ;
   RECT 0.00 275.31 179.36 277.02 ;
   RECT 0.00 277.02 179.36 278.73 ;
   RECT 0.00 278.73 179.36 280.44 ;
   RECT 0.00 280.44 179.36 282.15 ;
   RECT 0.00 282.15 179.36 283.86 ;
   RECT 0.00 283.86 179.36 285.57 ;
   RECT 0.00 285.57 179.36 287.28 ;
   RECT 0.00 287.28 179.36 288.99 ;
   RECT 0.00 288.99 179.36 290.70 ;
   RECT 0.00 290.70 179.36 292.41 ;
   RECT 0.00 292.41 179.36 294.12 ;
   RECT 0.00 294.12 179.36 295.83 ;
   RECT 0.00 295.83 179.36 297.54 ;
   RECT 0.00 297.54 179.36 299.25 ;
   RECT 0.00 299.25 179.36 300.96 ;
   RECT 0.00 300.96 179.36 302.67 ;
   RECT 0.00 302.67 179.36 304.38 ;
   RECT 0.00 304.38 179.36 306.09 ;
   RECT 0.00 306.09 179.36 307.80 ;
   RECT 0.00 307.80 179.36 309.51 ;
   RECT 0.00 309.51 179.36 311.22 ;
   RECT 0.00 311.22 179.36 312.93 ;
   RECT 0.00 312.93 179.36 314.64 ;
   RECT 0.00 314.64 179.36 316.35 ;
   RECT 0.00 316.35 179.36 318.06 ;
   RECT 0.00 318.06 179.36 319.77 ;
   RECT 0.00 319.77 179.36 321.48 ;
   RECT 0.00 321.48 179.36 323.19 ;
   RECT 0.00 323.19 179.36 324.90 ;
   RECT 0.00 324.90 179.36 326.61 ;
   RECT 0.00 326.61 179.36 328.32 ;
   RECT 0.00 328.32 179.36 330.03 ;
   RECT 0.00 330.03 179.36 331.74 ;
   RECT 0.00 331.74 179.36 333.45 ;
   RECT 0.00 333.45 179.36 335.16 ;
   RECT 0.00 335.16 179.36 336.87 ;
   RECT 0.00 336.87 179.36 338.58 ;
   RECT 0.00 338.58 179.36 340.29 ;
   RECT 0.00 340.29 179.36 342.00 ;
   RECT 0.00 342.00 179.36 343.71 ;
   RECT 0.00 343.71 179.36 345.42 ;
   RECT 0.00 345.42 179.36 347.13 ;
   RECT 0.00 347.13 179.36 348.84 ;
   RECT 0.00 348.84 179.36 350.55 ;
   RECT 0.00 350.55 179.36 352.26 ;
   RECT 0.00 352.26 179.36 353.97 ;
   RECT 0.00 353.97 179.36 355.68 ;
   RECT 0.00 355.68 179.36 357.39 ;
   RECT 0.00 357.39 179.36 359.10 ;
   RECT 0.00 359.10 179.36 360.81 ;
   RECT 0.00 360.81 179.36 362.52 ;
   RECT 0.00 362.52 179.36 364.23 ;
   RECT 0.00 364.23 179.36 365.94 ;
   RECT 0.00 365.94 179.36 367.65 ;
   RECT 0.00 367.65 179.36 369.36 ;
   RECT 0.00 369.36 179.36 371.07 ;
   RECT 0.00 371.07 179.36 372.78 ;
   RECT 0.00 372.78 179.36 374.49 ;
   RECT 0.00 374.49 179.36 376.20 ;
   RECT 0.00 376.20 179.36 377.91 ;
   RECT 0.00 377.91 179.36 379.62 ;
   RECT 0.00 379.62 179.36 381.33 ;
   RECT 0.00 381.33 179.36 383.04 ;
   RECT 0.00 383.04 179.36 384.75 ;
   RECT 0.00 384.75 179.36 386.46 ;
   RECT 0.00 386.46 179.36 388.17 ;
   RECT 0.00 388.17 179.36 389.88 ;
   RECT 0.00 389.88 179.36 391.59 ;
   RECT 0.00 391.59 179.36 393.30 ;
   RECT 0.00 393.30 179.36 395.01 ;
   RECT 0.00 395.01 179.36 396.72 ;
   RECT 0.00 396.72 179.36 398.43 ;
   RECT 0.00 398.43 179.36 400.14 ;
   RECT 0.00 400.14 179.36 401.85 ;
   RECT 0.00 401.85 202.54 403.56 ;
   RECT 0.00 403.56 202.54 405.27 ;
   RECT 0.00 405.27 202.54 406.98 ;
   RECT 0.00 406.98 202.54 408.69 ;
   RECT 0.00 408.69 202.54 410.40 ;
   RECT 0.00 410.40 202.54 412.11 ;
   RECT 0.00 412.11 202.54 413.82 ;
   RECT 0.00 413.82 202.54 415.53 ;
   RECT 0.00 415.53 202.54 417.24 ;
   RECT 0.00 417.24 202.54 418.95 ;
   RECT 0.00 418.95 202.54 420.66 ;
   RECT 0.00 420.66 202.54 422.37 ;
   RECT 0.00 422.37 202.54 424.08 ;
   RECT 0.00 424.08 202.54 425.79 ;
   RECT 0.00 425.79 202.54 427.50 ;
   RECT 0.00 427.50 202.54 429.21 ;
   RECT 0.00 429.21 202.54 430.92 ;
   RECT 0.00 430.92 179.36 432.63 ;
   RECT 0.00 432.63 179.36 434.34 ;
   RECT 0.00 434.34 179.36 436.05 ;
   RECT 0.00 436.05 179.36 437.76 ;
   RECT 0.00 437.76 179.36 439.47 ;
   RECT 0.00 439.47 179.36 441.18 ;
   RECT 0.00 441.18 179.36 442.89 ;
   RECT 0.00 442.89 179.36 444.60 ;
   RECT 0.00 444.60 179.36 446.31 ;
   RECT 0.00 446.31 179.36 448.02 ;
   RECT 0.00 448.02 179.36 449.73 ;
   RECT 0.00 449.73 179.36 451.44 ;
   RECT 0.00 451.44 179.36 453.15 ;
   RECT 0.00 453.15 179.36 454.86 ;
   RECT 0.00 454.86 179.36 456.57 ;
   RECT 0.00 456.57 179.36 458.28 ;
   RECT 0.00 458.28 179.36 459.99 ;
   RECT 0.00 459.99 179.36 461.70 ;
   RECT 0.00 461.70 179.36 463.41 ;
   RECT 0.00 463.41 179.36 465.12 ;
   RECT 0.00 465.12 179.36 466.83 ;
   RECT 0.00 466.83 179.36 468.54 ;
   RECT 0.00 468.54 179.36 470.25 ;
   RECT 0.00 470.25 179.36 471.96 ;
   RECT 0.00 471.96 179.36 473.67 ;
   RECT 0.00 473.67 179.36 475.38 ;
   RECT 0.00 475.38 179.36 477.09 ;
   RECT 0.00 477.09 179.36 478.80 ;
   RECT 0.00 478.80 179.36 480.51 ;
   RECT 0.00 480.51 179.36 482.22 ;
   RECT 0.00 482.22 179.36 483.93 ;
   RECT 0.00 483.93 179.36 485.64 ;
   RECT 0.00 485.64 179.36 487.35 ;
   RECT 0.00 487.35 179.36 489.06 ;
   RECT 0.00 489.06 179.36 490.77 ;
   RECT 0.00 490.77 179.36 492.48 ;
   RECT 0.00 492.48 179.36 494.19 ;
   RECT 0.00 494.19 179.36 495.90 ;
   RECT 0.00 495.90 179.36 497.61 ;
   RECT 0.00 497.61 179.36 499.32 ;
   RECT 0.00 499.32 179.36 501.03 ;
   RECT 0.00 501.03 179.36 502.74 ;
   RECT 0.00 502.74 179.36 504.45 ;
   RECT 0.00 504.45 179.36 506.16 ;
   RECT 0.00 506.16 179.36 507.87 ;
   RECT 0.00 507.87 179.36 509.58 ;
   RECT 0.00 509.58 179.36 511.29 ;
   RECT 0.00 511.29 179.36 513.00 ;
   RECT 0.00 513.00 179.36 514.71 ;
   RECT 0.00 514.71 179.36 516.42 ;
   RECT 0.00 516.42 179.36 518.13 ;
   RECT 0.00 518.13 179.36 519.84 ;
   RECT 0.00 519.84 179.36 521.55 ;
   RECT 0.00 521.55 179.36 523.26 ;
   RECT 0.00 523.26 179.36 524.97 ;
   RECT 0.00 524.97 179.36 526.68 ;
   RECT 0.00 526.68 179.36 528.39 ;
   RECT 0.00 528.39 179.36 530.10 ;
   RECT 0.00 530.10 179.36 531.81 ;
   RECT 0.00 531.81 179.36 533.52 ;
   RECT 0.00 533.52 179.36 535.23 ;
   RECT 0.00 535.23 179.36 536.94 ;
   RECT 0.00 536.94 179.36 538.65 ;
   RECT 0.00 538.65 179.36 540.36 ;
   RECT 0.00 540.36 179.36 542.07 ;
   RECT 0.00 542.07 179.36 543.78 ;
   RECT 0.00 543.78 179.36 545.49 ;
   RECT 0.00 545.49 179.36 547.20 ;
   RECT 0.00 547.20 179.36 548.91 ;
   RECT 0.00 548.91 179.36 550.62 ;
   RECT 0.00 550.62 179.36 552.33 ;
   RECT 0.00 552.33 179.36 554.04 ;
   RECT 0.00 554.04 179.36 555.75 ;
   RECT 0.00 555.75 179.36 557.46 ;
   RECT 0.00 557.46 179.36 559.17 ;
   RECT 0.00 559.17 179.36 560.88 ;
   RECT 0.00 560.88 179.36 562.59 ;
   RECT 0.00 562.59 179.36 564.30 ;
   RECT 0.00 564.30 179.36 566.01 ;
   RECT 0.00 566.01 179.36 567.72 ;
   RECT 0.00 567.72 179.36 569.43 ;
   RECT 0.00 569.43 179.36 571.14 ;
   RECT 0.00 571.14 179.36 572.85 ;
   RECT 0.00 572.85 179.36 574.56 ;
   RECT 0.00 574.56 179.36 576.27 ;
   RECT 0.00 576.27 179.36 577.98 ;
   RECT 0.00 577.98 179.36 579.69 ;
   RECT 0.00 579.69 179.36 581.40 ;
   RECT 0.00 581.40 179.36 583.11 ;
   RECT 0.00 583.11 179.36 584.82 ;
   RECT 0.00 584.82 179.36 586.53 ;
   RECT 0.00 586.53 179.36 588.24 ;
   RECT 0.00 588.24 179.36 589.95 ;
   RECT 0.00 589.95 179.36 591.66 ;
   RECT 0.00 591.66 179.36 593.37 ;
   RECT 0.00 593.37 179.36 595.08 ;
   RECT 0.00 595.08 179.36 596.79 ;
   RECT 0.00 596.79 179.36 598.50 ;
   RECT 0.00 598.50 179.36 600.21 ;
   RECT 0.00 600.21 179.36 601.92 ;
   RECT 0.00 601.92 179.36 603.63 ;
   RECT 0.00 603.63 179.36 605.34 ;
   RECT 0.00 605.34 179.36 607.05 ;
   RECT 0.00 607.05 179.36 608.76 ;
   RECT 0.00 608.76 179.36 610.47 ;
   RECT 0.00 610.47 179.36 612.18 ;
   RECT 0.00 612.18 179.36 613.89 ;
   RECT 0.00 613.89 179.36 615.60 ;
   RECT 0.00 615.60 179.36 617.31 ;
   RECT 0.00 617.31 179.36 619.02 ;
   RECT 0.00 619.02 179.36 620.73 ;
   RECT 0.00 620.73 179.36 622.44 ;
   RECT 0.00 622.44 179.36 624.15 ;
   RECT 0.00 624.15 179.36 625.86 ;
   RECT 0.00 625.86 179.36 627.57 ;
   RECT 0.00 627.57 179.36 629.28 ;
   RECT 0.00 629.28 179.36 630.99 ;
   RECT 0.00 630.99 179.36 632.70 ;
   RECT 0.00 632.70 179.36 634.41 ;
   RECT 0.00 634.41 179.36 636.12 ;
   RECT 0.00 636.12 179.36 637.83 ;
   RECT 0.00 637.83 179.36 639.54 ;
   RECT 0.00 639.54 179.36 641.25 ;
   RECT 0.00 641.25 179.36 642.96 ;
   RECT 0.00 642.96 179.36 644.67 ;
   RECT 0.00 644.67 179.36 646.38 ;
   RECT 0.00 646.38 179.36 648.09 ;
   RECT 0.00 648.09 179.36 649.80 ;
   RECT 0.00 649.80 179.36 651.51 ;
   RECT 0.00 651.51 179.36 653.22 ;
   RECT 0.00 653.22 179.36 654.93 ;
   RECT 0.00 654.93 179.36 656.64 ;
   RECT 0.00 656.64 179.36 658.35 ;
   RECT 0.00 658.35 179.36 660.06 ;
   RECT 0.00 660.06 179.36 661.77 ;
   RECT 0.00 661.77 179.36 663.48 ;
   RECT 0.00 663.48 179.36 665.19 ;
   RECT 0.00 665.19 179.36 666.90 ;
   RECT 0.00 666.90 179.36 668.61 ;
   RECT 0.00 668.61 179.36 670.32 ;
   RECT 0.00 670.32 179.36 672.03 ;
   RECT 0.00 672.03 179.36 673.74 ;
   RECT 0.00 673.74 179.36 675.45 ;
   RECT 0.00 675.45 179.36 677.16 ;
   RECT 0.00 677.16 179.36 678.87 ;
   RECT 0.00 678.87 179.36 680.58 ;
   RECT 0.00 680.58 179.36 682.29 ;
   RECT 0.00 682.29 179.36 684.00 ;
   RECT 0.00 684.00 179.36 685.71 ;
   RECT 0.00 685.71 179.36 687.42 ;
   RECT 0.00 687.42 179.36 689.13 ;
   RECT 0.00 689.13 179.36 690.84 ;
   RECT 0.00 690.84 179.36 692.55 ;
   RECT 0.00 692.55 179.36 694.26 ;
   RECT 0.00 694.26 179.36 695.97 ;
   RECT 0.00 695.97 179.36 697.68 ;
   RECT 0.00 697.68 179.36 699.39 ;
   RECT 0.00 699.39 179.36 701.10 ;
   RECT 0.00 701.10 179.36 702.81 ;
   RECT 0.00 702.81 179.36 704.52 ;
   RECT 0.00 704.52 179.36 706.23 ;
   RECT 0.00 706.23 179.36 707.94 ;
   RECT 0.00 707.94 179.36 709.65 ;
   RECT 0.00 709.65 179.36 711.36 ;
   RECT 0.00 711.36 179.36 713.07 ;
   RECT 0.00 713.07 179.36 714.78 ;
   RECT 0.00 714.78 179.36 716.49 ;
   RECT 0.00 716.49 179.36 718.20 ;
   RECT 0.00 718.20 179.36 719.91 ;
   RECT 0.00 719.91 179.36 721.62 ;
   RECT 0.00 721.62 179.36 723.33 ;
   RECT 0.00 723.33 179.36 725.04 ;
   RECT 0.00 725.04 179.36 726.75 ;
   RECT 0.00 726.75 179.36 728.46 ;
   RECT 0.00 728.46 179.36 730.17 ;
   RECT 0.00 730.17 179.36 731.88 ;
   RECT 0.00 731.88 179.36 733.59 ;
   RECT 0.00 733.59 179.36 735.30 ;
   RECT 0.00 735.30 179.36 737.01 ;
   RECT 0.00 737.01 179.36 738.72 ;
   RECT 0.00 738.72 179.36 740.43 ;
   RECT 0.00 740.43 179.36 742.14 ;
   RECT 0.00 742.14 179.36 743.85 ;
   RECT 0.00 743.85 179.36 745.56 ;
   RECT 0.00 745.56 179.36 747.27 ;
   RECT 0.00 747.27 179.36 748.98 ;
   RECT 0.00 748.98 179.36 750.69 ;
   RECT 0.00 750.69 179.36 752.40 ;
   RECT 0.00 752.40 179.36 754.11 ;
   RECT 0.00 754.11 179.36 755.82 ;
   RECT 0.00 755.82 179.36 757.53 ;
   RECT 0.00 757.53 179.36 759.24 ;
   RECT 0.00 759.24 179.36 760.95 ;
   RECT 0.00 760.95 179.36 762.66 ;
   RECT 0.00 762.66 179.36 764.37 ;
   RECT 0.00 764.37 179.36 766.08 ;
   RECT 0.00 766.08 179.36 767.79 ;
   RECT 0.00 767.79 179.36 769.50 ;
   RECT 0.00 769.50 179.36 771.21 ;
   RECT 0.00 771.21 179.36 772.92 ;
   RECT 0.00 772.92 179.36 774.63 ;
   RECT 0.00 774.63 179.36 776.34 ;
   RECT 0.00 776.34 179.36 778.05 ;
   RECT 0.00 778.05 179.36 779.76 ;
   RECT 0.00 779.76 179.36 781.47 ;
   RECT 0.00 781.47 179.36 783.18 ;
   RECT 0.00 783.18 179.36 784.89 ;
   RECT 0.00 784.89 179.36 786.60 ;
   RECT 0.00 786.60 179.36 788.31 ;
   RECT 0.00 788.31 179.36 790.02 ;
   RECT 0.00 790.02 179.36 791.73 ;
   RECT 0.00 791.73 179.36 793.44 ;
   RECT 0.00 793.44 179.36 795.15 ;
   RECT 0.00 795.15 179.36 796.86 ;
   RECT 0.00 796.86 179.36 798.57 ;
   RECT 0.00 798.57 179.36 800.28 ;
   RECT 0.00 800.28 179.36 801.99 ;
   RECT 0.00 801.99 179.36 803.70 ;
   RECT 0.00 803.70 179.36 805.41 ;
   RECT 0.00 805.41 179.36 807.12 ;
   RECT 0.00 807.12 179.36 808.83 ;
   RECT 0.00 808.83 179.36 810.54 ;
   RECT 0.00 810.54 179.36 812.25 ;
   RECT 0.00 812.25 179.36 813.96 ;
   RECT 0.00 813.96 179.36 815.67 ;
   RECT 0.00 815.67 179.36 817.38 ;
   RECT 0.00 817.38 179.36 819.09 ;
   RECT 0.00 819.09 179.36 820.80 ;
   RECT 0.00 820.80 179.36 822.51 ;
   RECT 0.00 822.51 179.36 824.22 ;
   RECT 0.00 824.22 179.36 825.93 ;
   RECT 0.00 825.93 179.36 827.64 ;
   RECT 0.00 827.64 179.36 829.35 ;
   RECT 0.00 829.35 179.36 831.06 ;
   RECT 0.00 831.06 179.36 832.77 ;
   RECT 0.00 832.77 179.36 834.48 ;
   RECT 0.00 834.48 179.36 836.19 ;
   RECT 0.00 836.19 179.36 837.90 ;
   RECT 0.00 837.90 179.36 839.61 ;
   RECT 0.00 839.61 179.36 841.32 ;
  LAYER via3 ;
   RECT 0.00 0.00 179.36 1.71 ;
   RECT 0.00 1.71 179.36 3.42 ;
   RECT 0.00 3.42 179.36 5.13 ;
   RECT 0.00 5.13 179.36 6.84 ;
   RECT 0.00 6.84 179.36 8.55 ;
   RECT 0.00 8.55 179.36 10.26 ;
   RECT 0.00 10.26 179.36 11.97 ;
   RECT 0.00 11.97 179.36 13.68 ;
   RECT 0.00 13.68 179.36 15.39 ;
   RECT 0.00 15.39 179.36 17.10 ;
   RECT 0.00 17.10 179.36 18.81 ;
   RECT 0.00 18.81 179.36 20.52 ;
   RECT 0.00 20.52 179.36 22.23 ;
   RECT 0.00 22.23 179.36 23.94 ;
   RECT 0.00 23.94 179.36 25.65 ;
   RECT 0.00 25.65 179.36 27.36 ;
   RECT 0.00 27.36 179.36 29.07 ;
   RECT 0.00 29.07 179.36 30.78 ;
   RECT 0.00 30.78 179.36 32.49 ;
   RECT 0.00 32.49 179.36 34.20 ;
   RECT 0.00 34.20 179.36 35.91 ;
   RECT 0.00 35.91 179.36 37.62 ;
   RECT 0.00 37.62 179.36 39.33 ;
   RECT 0.00 39.33 179.36 41.04 ;
   RECT 0.00 41.04 179.36 42.75 ;
   RECT 0.00 42.75 179.36 44.46 ;
   RECT 0.00 44.46 179.36 46.17 ;
   RECT 0.00 46.17 179.36 47.88 ;
   RECT 0.00 47.88 179.36 49.59 ;
   RECT 0.00 49.59 179.36 51.30 ;
   RECT 0.00 51.30 179.36 53.01 ;
   RECT 0.00 53.01 179.36 54.72 ;
   RECT 0.00 54.72 179.36 56.43 ;
   RECT 0.00 56.43 179.36 58.14 ;
   RECT 0.00 58.14 179.36 59.85 ;
   RECT 0.00 59.85 179.36 61.56 ;
   RECT 0.00 61.56 179.36 63.27 ;
   RECT 0.00 63.27 179.36 64.98 ;
   RECT 0.00 64.98 179.36 66.69 ;
   RECT 0.00 66.69 179.36 68.40 ;
   RECT 0.00 68.40 179.36 70.11 ;
   RECT 0.00 70.11 179.36 71.82 ;
   RECT 0.00 71.82 179.36 73.53 ;
   RECT 0.00 73.53 179.36 75.24 ;
   RECT 0.00 75.24 179.36 76.95 ;
   RECT 0.00 76.95 179.36 78.66 ;
   RECT 0.00 78.66 179.36 80.37 ;
   RECT 0.00 80.37 179.36 82.08 ;
   RECT 0.00 82.08 179.36 83.79 ;
   RECT 0.00 83.79 179.36 85.50 ;
   RECT 0.00 85.50 179.36 87.21 ;
   RECT 0.00 87.21 179.36 88.92 ;
   RECT 0.00 88.92 179.36 90.63 ;
   RECT 0.00 90.63 179.36 92.34 ;
   RECT 0.00 92.34 179.36 94.05 ;
   RECT 0.00 94.05 179.36 95.76 ;
   RECT 0.00 95.76 179.36 97.47 ;
   RECT 0.00 97.47 179.36 99.18 ;
   RECT 0.00 99.18 179.36 100.89 ;
   RECT 0.00 100.89 179.36 102.60 ;
   RECT 0.00 102.60 179.36 104.31 ;
   RECT 0.00 104.31 179.36 106.02 ;
   RECT 0.00 106.02 179.36 107.73 ;
   RECT 0.00 107.73 179.36 109.44 ;
   RECT 0.00 109.44 179.36 111.15 ;
   RECT 0.00 111.15 179.36 112.86 ;
   RECT 0.00 112.86 179.36 114.57 ;
   RECT 0.00 114.57 179.36 116.28 ;
   RECT 0.00 116.28 179.36 117.99 ;
   RECT 0.00 117.99 179.36 119.70 ;
   RECT 0.00 119.70 179.36 121.41 ;
   RECT 0.00 121.41 179.36 123.12 ;
   RECT 0.00 123.12 179.36 124.83 ;
   RECT 0.00 124.83 179.36 126.54 ;
   RECT 0.00 126.54 179.36 128.25 ;
   RECT 0.00 128.25 179.36 129.96 ;
   RECT 0.00 129.96 179.36 131.67 ;
   RECT 0.00 131.67 179.36 133.38 ;
   RECT 0.00 133.38 179.36 135.09 ;
   RECT 0.00 135.09 179.36 136.80 ;
   RECT 0.00 136.80 179.36 138.51 ;
   RECT 0.00 138.51 179.36 140.22 ;
   RECT 0.00 140.22 179.36 141.93 ;
   RECT 0.00 141.93 179.36 143.64 ;
   RECT 0.00 143.64 179.36 145.35 ;
   RECT 0.00 145.35 179.36 147.06 ;
   RECT 0.00 147.06 179.36 148.77 ;
   RECT 0.00 148.77 179.36 150.48 ;
   RECT 0.00 150.48 179.36 152.19 ;
   RECT 0.00 152.19 179.36 153.90 ;
   RECT 0.00 153.90 179.36 155.61 ;
   RECT 0.00 155.61 179.36 157.32 ;
   RECT 0.00 157.32 179.36 159.03 ;
   RECT 0.00 159.03 179.36 160.74 ;
   RECT 0.00 160.74 179.36 162.45 ;
   RECT 0.00 162.45 179.36 164.16 ;
   RECT 0.00 164.16 179.36 165.87 ;
   RECT 0.00 165.87 179.36 167.58 ;
   RECT 0.00 167.58 179.36 169.29 ;
   RECT 0.00 169.29 179.36 171.00 ;
   RECT 0.00 171.00 179.36 172.71 ;
   RECT 0.00 172.71 179.36 174.42 ;
   RECT 0.00 174.42 179.36 176.13 ;
   RECT 0.00 176.13 179.36 177.84 ;
   RECT 0.00 177.84 179.36 179.55 ;
   RECT 0.00 179.55 179.36 181.26 ;
   RECT 0.00 181.26 179.36 182.97 ;
   RECT 0.00 182.97 179.36 184.68 ;
   RECT 0.00 184.68 179.36 186.39 ;
   RECT 0.00 186.39 179.36 188.10 ;
   RECT 0.00 188.10 179.36 189.81 ;
   RECT 0.00 189.81 179.36 191.52 ;
   RECT 0.00 191.52 179.36 193.23 ;
   RECT 0.00 193.23 179.36 194.94 ;
   RECT 0.00 194.94 179.36 196.65 ;
   RECT 0.00 196.65 179.36 198.36 ;
   RECT 0.00 198.36 179.36 200.07 ;
   RECT 0.00 200.07 179.36 201.78 ;
   RECT 0.00 201.78 179.36 203.49 ;
   RECT 0.00 203.49 179.36 205.20 ;
   RECT 0.00 205.20 179.36 206.91 ;
   RECT 0.00 206.91 179.36 208.62 ;
   RECT 0.00 208.62 179.36 210.33 ;
   RECT 0.00 210.33 179.36 212.04 ;
   RECT 0.00 212.04 179.36 213.75 ;
   RECT 0.00 213.75 179.36 215.46 ;
   RECT 0.00 215.46 179.36 217.17 ;
   RECT 0.00 217.17 179.36 218.88 ;
   RECT 0.00 218.88 179.36 220.59 ;
   RECT 0.00 220.59 179.36 222.30 ;
   RECT 0.00 222.30 179.36 224.01 ;
   RECT 0.00 224.01 179.36 225.72 ;
   RECT 0.00 225.72 179.36 227.43 ;
   RECT 0.00 227.43 179.36 229.14 ;
   RECT 0.00 229.14 179.36 230.85 ;
   RECT 0.00 230.85 179.36 232.56 ;
   RECT 0.00 232.56 179.36 234.27 ;
   RECT 0.00 234.27 179.36 235.98 ;
   RECT 0.00 235.98 179.36 237.69 ;
   RECT 0.00 237.69 179.36 239.40 ;
   RECT 0.00 239.40 179.36 241.11 ;
   RECT 0.00 241.11 179.36 242.82 ;
   RECT 0.00 242.82 179.36 244.53 ;
   RECT 0.00 244.53 179.36 246.24 ;
   RECT 0.00 246.24 179.36 247.95 ;
   RECT 0.00 247.95 179.36 249.66 ;
   RECT 0.00 249.66 179.36 251.37 ;
   RECT 0.00 251.37 179.36 253.08 ;
   RECT 0.00 253.08 179.36 254.79 ;
   RECT 0.00 254.79 179.36 256.50 ;
   RECT 0.00 256.50 179.36 258.21 ;
   RECT 0.00 258.21 179.36 259.92 ;
   RECT 0.00 259.92 179.36 261.63 ;
   RECT 0.00 261.63 179.36 263.34 ;
   RECT 0.00 263.34 179.36 265.05 ;
   RECT 0.00 265.05 179.36 266.76 ;
   RECT 0.00 266.76 179.36 268.47 ;
   RECT 0.00 268.47 179.36 270.18 ;
   RECT 0.00 270.18 179.36 271.89 ;
   RECT 0.00 271.89 179.36 273.60 ;
   RECT 0.00 273.60 179.36 275.31 ;
   RECT 0.00 275.31 179.36 277.02 ;
   RECT 0.00 277.02 179.36 278.73 ;
   RECT 0.00 278.73 179.36 280.44 ;
   RECT 0.00 280.44 179.36 282.15 ;
   RECT 0.00 282.15 179.36 283.86 ;
   RECT 0.00 283.86 179.36 285.57 ;
   RECT 0.00 285.57 179.36 287.28 ;
   RECT 0.00 287.28 179.36 288.99 ;
   RECT 0.00 288.99 179.36 290.70 ;
   RECT 0.00 290.70 179.36 292.41 ;
   RECT 0.00 292.41 179.36 294.12 ;
   RECT 0.00 294.12 179.36 295.83 ;
   RECT 0.00 295.83 179.36 297.54 ;
   RECT 0.00 297.54 179.36 299.25 ;
   RECT 0.00 299.25 179.36 300.96 ;
   RECT 0.00 300.96 179.36 302.67 ;
   RECT 0.00 302.67 179.36 304.38 ;
   RECT 0.00 304.38 179.36 306.09 ;
   RECT 0.00 306.09 179.36 307.80 ;
   RECT 0.00 307.80 179.36 309.51 ;
   RECT 0.00 309.51 179.36 311.22 ;
   RECT 0.00 311.22 179.36 312.93 ;
   RECT 0.00 312.93 179.36 314.64 ;
   RECT 0.00 314.64 179.36 316.35 ;
   RECT 0.00 316.35 179.36 318.06 ;
   RECT 0.00 318.06 179.36 319.77 ;
   RECT 0.00 319.77 179.36 321.48 ;
   RECT 0.00 321.48 179.36 323.19 ;
   RECT 0.00 323.19 179.36 324.90 ;
   RECT 0.00 324.90 179.36 326.61 ;
   RECT 0.00 326.61 179.36 328.32 ;
   RECT 0.00 328.32 179.36 330.03 ;
   RECT 0.00 330.03 179.36 331.74 ;
   RECT 0.00 331.74 179.36 333.45 ;
   RECT 0.00 333.45 179.36 335.16 ;
   RECT 0.00 335.16 179.36 336.87 ;
   RECT 0.00 336.87 179.36 338.58 ;
   RECT 0.00 338.58 179.36 340.29 ;
   RECT 0.00 340.29 179.36 342.00 ;
   RECT 0.00 342.00 179.36 343.71 ;
   RECT 0.00 343.71 179.36 345.42 ;
   RECT 0.00 345.42 179.36 347.13 ;
   RECT 0.00 347.13 179.36 348.84 ;
   RECT 0.00 348.84 179.36 350.55 ;
   RECT 0.00 350.55 179.36 352.26 ;
   RECT 0.00 352.26 179.36 353.97 ;
   RECT 0.00 353.97 179.36 355.68 ;
   RECT 0.00 355.68 179.36 357.39 ;
   RECT 0.00 357.39 179.36 359.10 ;
   RECT 0.00 359.10 179.36 360.81 ;
   RECT 0.00 360.81 179.36 362.52 ;
   RECT 0.00 362.52 179.36 364.23 ;
   RECT 0.00 364.23 179.36 365.94 ;
   RECT 0.00 365.94 179.36 367.65 ;
   RECT 0.00 367.65 179.36 369.36 ;
   RECT 0.00 369.36 179.36 371.07 ;
   RECT 0.00 371.07 179.36 372.78 ;
   RECT 0.00 372.78 179.36 374.49 ;
   RECT 0.00 374.49 179.36 376.20 ;
   RECT 0.00 376.20 179.36 377.91 ;
   RECT 0.00 377.91 179.36 379.62 ;
   RECT 0.00 379.62 179.36 381.33 ;
   RECT 0.00 381.33 179.36 383.04 ;
   RECT 0.00 383.04 179.36 384.75 ;
   RECT 0.00 384.75 179.36 386.46 ;
   RECT 0.00 386.46 179.36 388.17 ;
   RECT 0.00 388.17 179.36 389.88 ;
   RECT 0.00 389.88 179.36 391.59 ;
   RECT 0.00 391.59 179.36 393.30 ;
   RECT 0.00 393.30 179.36 395.01 ;
   RECT 0.00 395.01 179.36 396.72 ;
   RECT 0.00 396.72 179.36 398.43 ;
   RECT 0.00 398.43 179.36 400.14 ;
   RECT 0.00 400.14 179.36 401.85 ;
   RECT 0.00 401.85 202.54 403.56 ;
   RECT 0.00 403.56 202.54 405.27 ;
   RECT 0.00 405.27 202.54 406.98 ;
   RECT 0.00 406.98 202.54 408.69 ;
   RECT 0.00 408.69 202.54 410.40 ;
   RECT 0.00 410.40 202.54 412.11 ;
   RECT 0.00 412.11 202.54 413.82 ;
   RECT 0.00 413.82 202.54 415.53 ;
   RECT 0.00 415.53 202.54 417.24 ;
   RECT 0.00 417.24 202.54 418.95 ;
   RECT 0.00 418.95 202.54 420.66 ;
   RECT 0.00 420.66 202.54 422.37 ;
   RECT 0.00 422.37 202.54 424.08 ;
   RECT 0.00 424.08 202.54 425.79 ;
   RECT 0.00 425.79 202.54 427.50 ;
   RECT 0.00 427.50 202.54 429.21 ;
   RECT 0.00 429.21 202.54 430.92 ;
   RECT 0.00 430.92 179.36 432.63 ;
   RECT 0.00 432.63 179.36 434.34 ;
   RECT 0.00 434.34 179.36 436.05 ;
   RECT 0.00 436.05 179.36 437.76 ;
   RECT 0.00 437.76 179.36 439.47 ;
   RECT 0.00 439.47 179.36 441.18 ;
   RECT 0.00 441.18 179.36 442.89 ;
   RECT 0.00 442.89 179.36 444.60 ;
   RECT 0.00 444.60 179.36 446.31 ;
   RECT 0.00 446.31 179.36 448.02 ;
   RECT 0.00 448.02 179.36 449.73 ;
   RECT 0.00 449.73 179.36 451.44 ;
   RECT 0.00 451.44 179.36 453.15 ;
   RECT 0.00 453.15 179.36 454.86 ;
   RECT 0.00 454.86 179.36 456.57 ;
   RECT 0.00 456.57 179.36 458.28 ;
   RECT 0.00 458.28 179.36 459.99 ;
   RECT 0.00 459.99 179.36 461.70 ;
   RECT 0.00 461.70 179.36 463.41 ;
   RECT 0.00 463.41 179.36 465.12 ;
   RECT 0.00 465.12 179.36 466.83 ;
   RECT 0.00 466.83 179.36 468.54 ;
   RECT 0.00 468.54 179.36 470.25 ;
   RECT 0.00 470.25 179.36 471.96 ;
   RECT 0.00 471.96 179.36 473.67 ;
   RECT 0.00 473.67 179.36 475.38 ;
   RECT 0.00 475.38 179.36 477.09 ;
   RECT 0.00 477.09 179.36 478.80 ;
   RECT 0.00 478.80 179.36 480.51 ;
   RECT 0.00 480.51 179.36 482.22 ;
   RECT 0.00 482.22 179.36 483.93 ;
   RECT 0.00 483.93 179.36 485.64 ;
   RECT 0.00 485.64 179.36 487.35 ;
   RECT 0.00 487.35 179.36 489.06 ;
   RECT 0.00 489.06 179.36 490.77 ;
   RECT 0.00 490.77 179.36 492.48 ;
   RECT 0.00 492.48 179.36 494.19 ;
   RECT 0.00 494.19 179.36 495.90 ;
   RECT 0.00 495.90 179.36 497.61 ;
   RECT 0.00 497.61 179.36 499.32 ;
   RECT 0.00 499.32 179.36 501.03 ;
   RECT 0.00 501.03 179.36 502.74 ;
   RECT 0.00 502.74 179.36 504.45 ;
   RECT 0.00 504.45 179.36 506.16 ;
   RECT 0.00 506.16 179.36 507.87 ;
   RECT 0.00 507.87 179.36 509.58 ;
   RECT 0.00 509.58 179.36 511.29 ;
   RECT 0.00 511.29 179.36 513.00 ;
   RECT 0.00 513.00 179.36 514.71 ;
   RECT 0.00 514.71 179.36 516.42 ;
   RECT 0.00 516.42 179.36 518.13 ;
   RECT 0.00 518.13 179.36 519.84 ;
   RECT 0.00 519.84 179.36 521.55 ;
   RECT 0.00 521.55 179.36 523.26 ;
   RECT 0.00 523.26 179.36 524.97 ;
   RECT 0.00 524.97 179.36 526.68 ;
   RECT 0.00 526.68 179.36 528.39 ;
   RECT 0.00 528.39 179.36 530.10 ;
   RECT 0.00 530.10 179.36 531.81 ;
   RECT 0.00 531.81 179.36 533.52 ;
   RECT 0.00 533.52 179.36 535.23 ;
   RECT 0.00 535.23 179.36 536.94 ;
   RECT 0.00 536.94 179.36 538.65 ;
   RECT 0.00 538.65 179.36 540.36 ;
   RECT 0.00 540.36 179.36 542.07 ;
   RECT 0.00 542.07 179.36 543.78 ;
   RECT 0.00 543.78 179.36 545.49 ;
   RECT 0.00 545.49 179.36 547.20 ;
   RECT 0.00 547.20 179.36 548.91 ;
   RECT 0.00 548.91 179.36 550.62 ;
   RECT 0.00 550.62 179.36 552.33 ;
   RECT 0.00 552.33 179.36 554.04 ;
   RECT 0.00 554.04 179.36 555.75 ;
   RECT 0.00 555.75 179.36 557.46 ;
   RECT 0.00 557.46 179.36 559.17 ;
   RECT 0.00 559.17 179.36 560.88 ;
   RECT 0.00 560.88 179.36 562.59 ;
   RECT 0.00 562.59 179.36 564.30 ;
   RECT 0.00 564.30 179.36 566.01 ;
   RECT 0.00 566.01 179.36 567.72 ;
   RECT 0.00 567.72 179.36 569.43 ;
   RECT 0.00 569.43 179.36 571.14 ;
   RECT 0.00 571.14 179.36 572.85 ;
   RECT 0.00 572.85 179.36 574.56 ;
   RECT 0.00 574.56 179.36 576.27 ;
   RECT 0.00 576.27 179.36 577.98 ;
   RECT 0.00 577.98 179.36 579.69 ;
   RECT 0.00 579.69 179.36 581.40 ;
   RECT 0.00 581.40 179.36 583.11 ;
   RECT 0.00 583.11 179.36 584.82 ;
   RECT 0.00 584.82 179.36 586.53 ;
   RECT 0.00 586.53 179.36 588.24 ;
   RECT 0.00 588.24 179.36 589.95 ;
   RECT 0.00 589.95 179.36 591.66 ;
   RECT 0.00 591.66 179.36 593.37 ;
   RECT 0.00 593.37 179.36 595.08 ;
   RECT 0.00 595.08 179.36 596.79 ;
   RECT 0.00 596.79 179.36 598.50 ;
   RECT 0.00 598.50 179.36 600.21 ;
   RECT 0.00 600.21 179.36 601.92 ;
   RECT 0.00 601.92 179.36 603.63 ;
   RECT 0.00 603.63 179.36 605.34 ;
   RECT 0.00 605.34 179.36 607.05 ;
   RECT 0.00 607.05 179.36 608.76 ;
   RECT 0.00 608.76 179.36 610.47 ;
   RECT 0.00 610.47 179.36 612.18 ;
   RECT 0.00 612.18 179.36 613.89 ;
   RECT 0.00 613.89 179.36 615.60 ;
   RECT 0.00 615.60 179.36 617.31 ;
   RECT 0.00 617.31 179.36 619.02 ;
   RECT 0.00 619.02 179.36 620.73 ;
   RECT 0.00 620.73 179.36 622.44 ;
   RECT 0.00 622.44 179.36 624.15 ;
   RECT 0.00 624.15 179.36 625.86 ;
   RECT 0.00 625.86 179.36 627.57 ;
   RECT 0.00 627.57 179.36 629.28 ;
   RECT 0.00 629.28 179.36 630.99 ;
   RECT 0.00 630.99 179.36 632.70 ;
   RECT 0.00 632.70 179.36 634.41 ;
   RECT 0.00 634.41 179.36 636.12 ;
   RECT 0.00 636.12 179.36 637.83 ;
   RECT 0.00 637.83 179.36 639.54 ;
   RECT 0.00 639.54 179.36 641.25 ;
   RECT 0.00 641.25 179.36 642.96 ;
   RECT 0.00 642.96 179.36 644.67 ;
   RECT 0.00 644.67 179.36 646.38 ;
   RECT 0.00 646.38 179.36 648.09 ;
   RECT 0.00 648.09 179.36 649.80 ;
   RECT 0.00 649.80 179.36 651.51 ;
   RECT 0.00 651.51 179.36 653.22 ;
   RECT 0.00 653.22 179.36 654.93 ;
   RECT 0.00 654.93 179.36 656.64 ;
   RECT 0.00 656.64 179.36 658.35 ;
   RECT 0.00 658.35 179.36 660.06 ;
   RECT 0.00 660.06 179.36 661.77 ;
   RECT 0.00 661.77 179.36 663.48 ;
   RECT 0.00 663.48 179.36 665.19 ;
   RECT 0.00 665.19 179.36 666.90 ;
   RECT 0.00 666.90 179.36 668.61 ;
   RECT 0.00 668.61 179.36 670.32 ;
   RECT 0.00 670.32 179.36 672.03 ;
   RECT 0.00 672.03 179.36 673.74 ;
   RECT 0.00 673.74 179.36 675.45 ;
   RECT 0.00 675.45 179.36 677.16 ;
   RECT 0.00 677.16 179.36 678.87 ;
   RECT 0.00 678.87 179.36 680.58 ;
   RECT 0.00 680.58 179.36 682.29 ;
   RECT 0.00 682.29 179.36 684.00 ;
   RECT 0.00 684.00 179.36 685.71 ;
   RECT 0.00 685.71 179.36 687.42 ;
   RECT 0.00 687.42 179.36 689.13 ;
   RECT 0.00 689.13 179.36 690.84 ;
   RECT 0.00 690.84 179.36 692.55 ;
   RECT 0.00 692.55 179.36 694.26 ;
   RECT 0.00 694.26 179.36 695.97 ;
   RECT 0.00 695.97 179.36 697.68 ;
   RECT 0.00 697.68 179.36 699.39 ;
   RECT 0.00 699.39 179.36 701.10 ;
   RECT 0.00 701.10 179.36 702.81 ;
   RECT 0.00 702.81 179.36 704.52 ;
   RECT 0.00 704.52 179.36 706.23 ;
   RECT 0.00 706.23 179.36 707.94 ;
   RECT 0.00 707.94 179.36 709.65 ;
   RECT 0.00 709.65 179.36 711.36 ;
   RECT 0.00 711.36 179.36 713.07 ;
   RECT 0.00 713.07 179.36 714.78 ;
   RECT 0.00 714.78 179.36 716.49 ;
   RECT 0.00 716.49 179.36 718.20 ;
   RECT 0.00 718.20 179.36 719.91 ;
   RECT 0.00 719.91 179.36 721.62 ;
   RECT 0.00 721.62 179.36 723.33 ;
   RECT 0.00 723.33 179.36 725.04 ;
   RECT 0.00 725.04 179.36 726.75 ;
   RECT 0.00 726.75 179.36 728.46 ;
   RECT 0.00 728.46 179.36 730.17 ;
   RECT 0.00 730.17 179.36 731.88 ;
   RECT 0.00 731.88 179.36 733.59 ;
   RECT 0.00 733.59 179.36 735.30 ;
   RECT 0.00 735.30 179.36 737.01 ;
   RECT 0.00 737.01 179.36 738.72 ;
   RECT 0.00 738.72 179.36 740.43 ;
   RECT 0.00 740.43 179.36 742.14 ;
   RECT 0.00 742.14 179.36 743.85 ;
   RECT 0.00 743.85 179.36 745.56 ;
   RECT 0.00 745.56 179.36 747.27 ;
   RECT 0.00 747.27 179.36 748.98 ;
   RECT 0.00 748.98 179.36 750.69 ;
   RECT 0.00 750.69 179.36 752.40 ;
   RECT 0.00 752.40 179.36 754.11 ;
   RECT 0.00 754.11 179.36 755.82 ;
   RECT 0.00 755.82 179.36 757.53 ;
   RECT 0.00 757.53 179.36 759.24 ;
   RECT 0.00 759.24 179.36 760.95 ;
   RECT 0.00 760.95 179.36 762.66 ;
   RECT 0.00 762.66 179.36 764.37 ;
   RECT 0.00 764.37 179.36 766.08 ;
   RECT 0.00 766.08 179.36 767.79 ;
   RECT 0.00 767.79 179.36 769.50 ;
   RECT 0.00 769.50 179.36 771.21 ;
   RECT 0.00 771.21 179.36 772.92 ;
   RECT 0.00 772.92 179.36 774.63 ;
   RECT 0.00 774.63 179.36 776.34 ;
   RECT 0.00 776.34 179.36 778.05 ;
   RECT 0.00 778.05 179.36 779.76 ;
   RECT 0.00 779.76 179.36 781.47 ;
   RECT 0.00 781.47 179.36 783.18 ;
   RECT 0.00 783.18 179.36 784.89 ;
   RECT 0.00 784.89 179.36 786.60 ;
   RECT 0.00 786.60 179.36 788.31 ;
   RECT 0.00 788.31 179.36 790.02 ;
   RECT 0.00 790.02 179.36 791.73 ;
   RECT 0.00 791.73 179.36 793.44 ;
   RECT 0.00 793.44 179.36 795.15 ;
   RECT 0.00 795.15 179.36 796.86 ;
   RECT 0.00 796.86 179.36 798.57 ;
   RECT 0.00 798.57 179.36 800.28 ;
   RECT 0.00 800.28 179.36 801.99 ;
   RECT 0.00 801.99 179.36 803.70 ;
   RECT 0.00 803.70 179.36 805.41 ;
   RECT 0.00 805.41 179.36 807.12 ;
   RECT 0.00 807.12 179.36 808.83 ;
   RECT 0.00 808.83 179.36 810.54 ;
   RECT 0.00 810.54 179.36 812.25 ;
   RECT 0.00 812.25 179.36 813.96 ;
   RECT 0.00 813.96 179.36 815.67 ;
   RECT 0.00 815.67 179.36 817.38 ;
   RECT 0.00 817.38 179.36 819.09 ;
   RECT 0.00 819.09 179.36 820.80 ;
   RECT 0.00 820.80 179.36 822.51 ;
   RECT 0.00 822.51 179.36 824.22 ;
   RECT 0.00 824.22 179.36 825.93 ;
   RECT 0.00 825.93 179.36 827.64 ;
   RECT 0.00 827.64 179.36 829.35 ;
   RECT 0.00 829.35 179.36 831.06 ;
   RECT 0.00 831.06 179.36 832.77 ;
   RECT 0.00 832.77 179.36 834.48 ;
   RECT 0.00 834.48 179.36 836.19 ;
   RECT 0.00 836.19 179.36 837.90 ;
   RECT 0.00 837.90 179.36 839.61 ;
   RECT 0.00 839.61 179.36 841.32 ;
  LAYER metal4 ;
   RECT 0.00 0.00 179.36 1.71 ;
   RECT 0.00 1.71 179.36 3.42 ;
   RECT 0.00 3.42 179.36 5.13 ;
   RECT 0.00 5.13 179.36 6.84 ;
   RECT 0.00 6.84 179.36 8.55 ;
   RECT 0.00 8.55 179.36 10.26 ;
   RECT 0.00 10.26 179.36 11.97 ;
   RECT 0.00 11.97 179.36 13.68 ;
   RECT 0.00 13.68 179.36 15.39 ;
   RECT 0.00 15.39 179.36 17.10 ;
   RECT 0.00 17.10 179.36 18.81 ;
   RECT 0.00 18.81 179.36 20.52 ;
   RECT 0.00 20.52 179.36 22.23 ;
   RECT 0.00 22.23 179.36 23.94 ;
   RECT 0.00 23.94 179.36 25.65 ;
   RECT 0.00 25.65 179.36 27.36 ;
   RECT 0.00 27.36 179.36 29.07 ;
   RECT 0.00 29.07 179.36 30.78 ;
   RECT 0.00 30.78 179.36 32.49 ;
   RECT 0.00 32.49 179.36 34.20 ;
   RECT 0.00 34.20 179.36 35.91 ;
   RECT 0.00 35.91 179.36 37.62 ;
   RECT 0.00 37.62 179.36 39.33 ;
   RECT 0.00 39.33 179.36 41.04 ;
   RECT 0.00 41.04 179.36 42.75 ;
   RECT 0.00 42.75 179.36 44.46 ;
   RECT 0.00 44.46 179.36 46.17 ;
   RECT 0.00 46.17 179.36 47.88 ;
   RECT 0.00 47.88 179.36 49.59 ;
   RECT 0.00 49.59 179.36 51.30 ;
   RECT 0.00 51.30 179.36 53.01 ;
   RECT 0.00 53.01 179.36 54.72 ;
   RECT 0.00 54.72 179.36 56.43 ;
   RECT 0.00 56.43 179.36 58.14 ;
   RECT 0.00 58.14 179.36 59.85 ;
   RECT 0.00 59.85 179.36 61.56 ;
   RECT 0.00 61.56 179.36 63.27 ;
   RECT 0.00 63.27 179.36 64.98 ;
   RECT 0.00 64.98 179.36 66.69 ;
   RECT 0.00 66.69 179.36 68.40 ;
   RECT 0.00 68.40 179.36 70.11 ;
   RECT 0.00 70.11 179.36 71.82 ;
   RECT 0.00 71.82 179.36 73.53 ;
   RECT 0.00 73.53 179.36 75.24 ;
   RECT 0.00 75.24 179.36 76.95 ;
   RECT 0.00 76.95 179.36 78.66 ;
   RECT 0.00 78.66 179.36 80.37 ;
   RECT 0.00 80.37 179.36 82.08 ;
   RECT 0.00 82.08 179.36 83.79 ;
   RECT 0.00 83.79 179.36 85.50 ;
   RECT 0.00 85.50 179.36 87.21 ;
   RECT 0.00 87.21 179.36 88.92 ;
   RECT 0.00 88.92 179.36 90.63 ;
   RECT 0.00 90.63 179.36 92.34 ;
   RECT 0.00 92.34 179.36 94.05 ;
   RECT 0.00 94.05 179.36 95.76 ;
   RECT 0.00 95.76 179.36 97.47 ;
   RECT 0.00 97.47 179.36 99.18 ;
   RECT 0.00 99.18 179.36 100.89 ;
   RECT 0.00 100.89 179.36 102.60 ;
   RECT 0.00 102.60 179.36 104.31 ;
   RECT 0.00 104.31 179.36 106.02 ;
   RECT 0.00 106.02 179.36 107.73 ;
   RECT 0.00 107.73 179.36 109.44 ;
   RECT 0.00 109.44 179.36 111.15 ;
   RECT 0.00 111.15 179.36 112.86 ;
   RECT 0.00 112.86 179.36 114.57 ;
   RECT 0.00 114.57 179.36 116.28 ;
   RECT 0.00 116.28 179.36 117.99 ;
   RECT 0.00 117.99 179.36 119.70 ;
   RECT 0.00 119.70 179.36 121.41 ;
   RECT 0.00 121.41 179.36 123.12 ;
   RECT 0.00 123.12 179.36 124.83 ;
   RECT 0.00 124.83 179.36 126.54 ;
   RECT 0.00 126.54 179.36 128.25 ;
   RECT 0.00 128.25 179.36 129.96 ;
   RECT 0.00 129.96 179.36 131.67 ;
   RECT 0.00 131.67 179.36 133.38 ;
   RECT 0.00 133.38 179.36 135.09 ;
   RECT 0.00 135.09 179.36 136.80 ;
   RECT 0.00 136.80 179.36 138.51 ;
   RECT 0.00 138.51 179.36 140.22 ;
   RECT 0.00 140.22 179.36 141.93 ;
   RECT 0.00 141.93 179.36 143.64 ;
   RECT 0.00 143.64 179.36 145.35 ;
   RECT 0.00 145.35 179.36 147.06 ;
   RECT 0.00 147.06 179.36 148.77 ;
   RECT 0.00 148.77 179.36 150.48 ;
   RECT 0.00 150.48 179.36 152.19 ;
   RECT 0.00 152.19 179.36 153.90 ;
   RECT 0.00 153.90 179.36 155.61 ;
   RECT 0.00 155.61 179.36 157.32 ;
   RECT 0.00 157.32 179.36 159.03 ;
   RECT 0.00 159.03 179.36 160.74 ;
   RECT 0.00 160.74 179.36 162.45 ;
   RECT 0.00 162.45 179.36 164.16 ;
   RECT 0.00 164.16 179.36 165.87 ;
   RECT 0.00 165.87 179.36 167.58 ;
   RECT 0.00 167.58 179.36 169.29 ;
   RECT 0.00 169.29 179.36 171.00 ;
   RECT 0.00 171.00 179.36 172.71 ;
   RECT 0.00 172.71 179.36 174.42 ;
   RECT 0.00 174.42 179.36 176.13 ;
   RECT 0.00 176.13 179.36 177.84 ;
   RECT 0.00 177.84 179.36 179.55 ;
   RECT 0.00 179.55 179.36 181.26 ;
   RECT 0.00 181.26 179.36 182.97 ;
   RECT 0.00 182.97 179.36 184.68 ;
   RECT 0.00 184.68 179.36 186.39 ;
   RECT 0.00 186.39 179.36 188.10 ;
   RECT 0.00 188.10 179.36 189.81 ;
   RECT 0.00 189.81 179.36 191.52 ;
   RECT 0.00 191.52 179.36 193.23 ;
   RECT 0.00 193.23 179.36 194.94 ;
   RECT 0.00 194.94 179.36 196.65 ;
   RECT 0.00 196.65 179.36 198.36 ;
   RECT 0.00 198.36 179.36 200.07 ;
   RECT 0.00 200.07 179.36 201.78 ;
   RECT 0.00 201.78 179.36 203.49 ;
   RECT 0.00 203.49 179.36 205.20 ;
   RECT 0.00 205.20 179.36 206.91 ;
   RECT 0.00 206.91 179.36 208.62 ;
   RECT 0.00 208.62 179.36 210.33 ;
   RECT 0.00 210.33 179.36 212.04 ;
   RECT 0.00 212.04 179.36 213.75 ;
   RECT 0.00 213.75 179.36 215.46 ;
   RECT 0.00 215.46 179.36 217.17 ;
   RECT 0.00 217.17 179.36 218.88 ;
   RECT 0.00 218.88 179.36 220.59 ;
   RECT 0.00 220.59 179.36 222.30 ;
   RECT 0.00 222.30 179.36 224.01 ;
   RECT 0.00 224.01 179.36 225.72 ;
   RECT 0.00 225.72 179.36 227.43 ;
   RECT 0.00 227.43 179.36 229.14 ;
   RECT 0.00 229.14 179.36 230.85 ;
   RECT 0.00 230.85 179.36 232.56 ;
   RECT 0.00 232.56 179.36 234.27 ;
   RECT 0.00 234.27 179.36 235.98 ;
   RECT 0.00 235.98 179.36 237.69 ;
   RECT 0.00 237.69 179.36 239.40 ;
   RECT 0.00 239.40 179.36 241.11 ;
   RECT 0.00 241.11 179.36 242.82 ;
   RECT 0.00 242.82 179.36 244.53 ;
   RECT 0.00 244.53 179.36 246.24 ;
   RECT 0.00 246.24 179.36 247.95 ;
   RECT 0.00 247.95 179.36 249.66 ;
   RECT 0.00 249.66 179.36 251.37 ;
   RECT 0.00 251.37 179.36 253.08 ;
   RECT 0.00 253.08 179.36 254.79 ;
   RECT 0.00 254.79 179.36 256.50 ;
   RECT 0.00 256.50 179.36 258.21 ;
   RECT 0.00 258.21 179.36 259.92 ;
   RECT 0.00 259.92 179.36 261.63 ;
   RECT 0.00 261.63 179.36 263.34 ;
   RECT 0.00 263.34 179.36 265.05 ;
   RECT 0.00 265.05 179.36 266.76 ;
   RECT 0.00 266.76 179.36 268.47 ;
   RECT 0.00 268.47 179.36 270.18 ;
   RECT 0.00 270.18 179.36 271.89 ;
   RECT 0.00 271.89 179.36 273.60 ;
   RECT 0.00 273.60 179.36 275.31 ;
   RECT 0.00 275.31 179.36 277.02 ;
   RECT 0.00 277.02 179.36 278.73 ;
   RECT 0.00 278.73 179.36 280.44 ;
   RECT 0.00 280.44 179.36 282.15 ;
   RECT 0.00 282.15 179.36 283.86 ;
   RECT 0.00 283.86 179.36 285.57 ;
   RECT 0.00 285.57 179.36 287.28 ;
   RECT 0.00 287.28 179.36 288.99 ;
   RECT 0.00 288.99 179.36 290.70 ;
   RECT 0.00 290.70 179.36 292.41 ;
   RECT 0.00 292.41 179.36 294.12 ;
   RECT 0.00 294.12 179.36 295.83 ;
   RECT 0.00 295.83 179.36 297.54 ;
   RECT 0.00 297.54 179.36 299.25 ;
   RECT 0.00 299.25 179.36 300.96 ;
   RECT 0.00 300.96 179.36 302.67 ;
   RECT 0.00 302.67 179.36 304.38 ;
   RECT 0.00 304.38 179.36 306.09 ;
   RECT 0.00 306.09 179.36 307.80 ;
   RECT 0.00 307.80 179.36 309.51 ;
   RECT 0.00 309.51 179.36 311.22 ;
   RECT 0.00 311.22 179.36 312.93 ;
   RECT 0.00 312.93 179.36 314.64 ;
   RECT 0.00 314.64 179.36 316.35 ;
   RECT 0.00 316.35 179.36 318.06 ;
   RECT 0.00 318.06 179.36 319.77 ;
   RECT 0.00 319.77 179.36 321.48 ;
   RECT 0.00 321.48 179.36 323.19 ;
   RECT 0.00 323.19 179.36 324.90 ;
   RECT 0.00 324.90 179.36 326.61 ;
   RECT 0.00 326.61 179.36 328.32 ;
   RECT 0.00 328.32 179.36 330.03 ;
   RECT 0.00 330.03 179.36 331.74 ;
   RECT 0.00 331.74 179.36 333.45 ;
   RECT 0.00 333.45 179.36 335.16 ;
   RECT 0.00 335.16 179.36 336.87 ;
   RECT 0.00 336.87 179.36 338.58 ;
   RECT 0.00 338.58 179.36 340.29 ;
   RECT 0.00 340.29 179.36 342.00 ;
   RECT 0.00 342.00 179.36 343.71 ;
   RECT 0.00 343.71 179.36 345.42 ;
   RECT 0.00 345.42 179.36 347.13 ;
   RECT 0.00 347.13 179.36 348.84 ;
   RECT 0.00 348.84 179.36 350.55 ;
   RECT 0.00 350.55 179.36 352.26 ;
   RECT 0.00 352.26 179.36 353.97 ;
   RECT 0.00 353.97 179.36 355.68 ;
   RECT 0.00 355.68 179.36 357.39 ;
   RECT 0.00 357.39 179.36 359.10 ;
   RECT 0.00 359.10 179.36 360.81 ;
   RECT 0.00 360.81 179.36 362.52 ;
   RECT 0.00 362.52 179.36 364.23 ;
   RECT 0.00 364.23 179.36 365.94 ;
   RECT 0.00 365.94 179.36 367.65 ;
   RECT 0.00 367.65 179.36 369.36 ;
   RECT 0.00 369.36 179.36 371.07 ;
   RECT 0.00 371.07 179.36 372.78 ;
   RECT 0.00 372.78 179.36 374.49 ;
   RECT 0.00 374.49 179.36 376.20 ;
   RECT 0.00 376.20 179.36 377.91 ;
   RECT 0.00 377.91 179.36 379.62 ;
   RECT 0.00 379.62 179.36 381.33 ;
   RECT 0.00 381.33 179.36 383.04 ;
   RECT 0.00 383.04 179.36 384.75 ;
   RECT 0.00 384.75 179.36 386.46 ;
   RECT 0.00 386.46 179.36 388.17 ;
   RECT 0.00 388.17 179.36 389.88 ;
   RECT 0.00 389.88 179.36 391.59 ;
   RECT 0.00 391.59 179.36 393.30 ;
   RECT 0.00 393.30 179.36 395.01 ;
   RECT 0.00 395.01 179.36 396.72 ;
   RECT 0.00 396.72 179.36 398.43 ;
   RECT 0.00 398.43 179.36 400.14 ;
   RECT 0.00 400.14 179.36 401.85 ;
   RECT 0.00 401.85 202.54 403.56 ;
   RECT 0.00 403.56 202.54 405.27 ;
   RECT 0.00 405.27 202.54 406.98 ;
   RECT 0.00 406.98 202.54 408.69 ;
   RECT 0.00 408.69 202.54 410.40 ;
   RECT 0.00 410.40 202.54 412.11 ;
   RECT 0.00 412.11 202.54 413.82 ;
   RECT 0.00 413.82 202.54 415.53 ;
   RECT 0.00 415.53 202.54 417.24 ;
   RECT 0.00 417.24 202.54 418.95 ;
   RECT 0.00 418.95 202.54 420.66 ;
   RECT 0.00 420.66 202.54 422.37 ;
   RECT 0.00 422.37 202.54 424.08 ;
   RECT 0.00 424.08 202.54 425.79 ;
   RECT 0.00 425.79 202.54 427.50 ;
   RECT 0.00 427.50 202.54 429.21 ;
   RECT 0.00 429.21 202.54 430.92 ;
   RECT 0.00 430.92 179.36 432.63 ;
   RECT 0.00 432.63 179.36 434.34 ;
   RECT 0.00 434.34 179.36 436.05 ;
   RECT 0.00 436.05 179.36 437.76 ;
   RECT 0.00 437.76 179.36 439.47 ;
   RECT 0.00 439.47 179.36 441.18 ;
   RECT 0.00 441.18 179.36 442.89 ;
   RECT 0.00 442.89 179.36 444.60 ;
   RECT 0.00 444.60 179.36 446.31 ;
   RECT 0.00 446.31 179.36 448.02 ;
   RECT 0.00 448.02 179.36 449.73 ;
   RECT 0.00 449.73 179.36 451.44 ;
   RECT 0.00 451.44 179.36 453.15 ;
   RECT 0.00 453.15 179.36 454.86 ;
   RECT 0.00 454.86 179.36 456.57 ;
   RECT 0.00 456.57 179.36 458.28 ;
   RECT 0.00 458.28 179.36 459.99 ;
   RECT 0.00 459.99 179.36 461.70 ;
   RECT 0.00 461.70 179.36 463.41 ;
   RECT 0.00 463.41 179.36 465.12 ;
   RECT 0.00 465.12 179.36 466.83 ;
   RECT 0.00 466.83 179.36 468.54 ;
   RECT 0.00 468.54 179.36 470.25 ;
   RECT 0.00 470.25 179.36 471.96 ;
   RECT 0.00 471.96 179.36 473.67 ;
   RECT 0.00 473.67 179.36 475.38 ;
   RECT 0.00 475.38 179.36 477.09 ;
   RECT 0.00 477.09 179.36 478.80 ;
   RECT 0.00 478.80 179.36 480.51 ;
   RECT 0.00 480.51 179.36 482.22 ;
   RECT 0.00 482.22 179.36 483.93 ;
   RECT 0.00 483.93 179.36 485.64 ;
   RECT 0.00 485.64 179.36 487.35 ;
   RECT 0.00 487.35 179.36 489.06 ;
   RECT 0.00 489.06 179.36 490.77 ;
   RECT 0.00 490.77 179.36 492.48 ;
   RECT 0.00 492.48 179.36 494.19 ;
   RECT 0.00 494.19 179.36 495.90 ;
   RECT 0.00 495.90 179.36 497.61 ;
   RECT 0.00 497.61 179.36 499.32 ;
   RECT 0.00 499.32 179.36 501.03 ;
   RECT 0.00 501.03 179.36 502.74 ;
   RECT 0.00 502.74 179.36 504.45 ;
   RECT 0.00 504.45 179.36 506.16 ;
   RECT 0.00 506.16 179.36 507.87 ;
   RECT 0.00 507.87 179.36 509.58 ;
   RECT 0.00 509.58 179.36 511.29 ;
   RECT 0.00 511.29 179.36 513.00 ;
   RECT 0.00 513.00 179.36 514.71 ;
   RECT 0.00 514.71 179.36 516.42 ;
   RECT 0.00 516.42 179.36 518.13 ;
   RECT 0.00 518.13 179.36 519.84 ;
   RECT 0.00 519.84 179.36 521.55 ;
   RECT 0.00 521.55 179.36 523.26 ;
   RECT 0.00 523.26 179.36 524.97 ;
   RECT 0.00 524.97 179.36 526.68 ;
   RECT 0.00 526.68 179.36 528.39 ;
   RECT 0.00 528.39 179.36 530.10 ;
   RECT 0.00 530.10 179.36 531.81 ;
   RECT 0.00 531.81 179.36 533.52 ;
   RECT 0.00 533.52 179.36 535.23 ;
   RECT 0.00 535.23 179.36 536.94 ;
   RECT 0.00 536.94 179.36 538.65 ;
   RECT 0.00 538.65 179.36 540.36 ;
   RECT 0.00 540.36 179.36 542.07 ;
   RECT 0.00 542.07 179.36 543.78 ;
   RECT 0.00 543.78 179.36 545.49 ;
   RECT 0.00 545.49 179.36 547.20 ;
   RECT 0.00 547.20 179.36 548.91 ;
   RECT 0.00 548.91 179.36 550.62 ;
   RECT 0.00 550.62 179.36 552.33 ;
   RECT 0.00 552.33 179.36 554.04 ;
   RECT 0.00 554.04 179.36 555.75 ;
   RECT 0.00 555.75 179.36 557.46 ;
   RECT 0.00 557.46 179.36 559.17 ;
   RECT 0.00 559.17 179.36 560.88 ;
   RECT 0.00 560.88 179.36 562.59 ;
   RECT 0.00 562.59 179.36 564.30 ;
   RECT 0.00 564.30 179.36 566.01 ;
   RECT 0.00 566.01 179.36 567.72 ;
   RECT 0.00 567.72 179.36 569.43 ;
   RECT 0.00 569.43 179.36 571.14 ;
   RECT 0.00 571.14 179.36 572.85 ;
   RECT 0.00 572.85 179.36 574.56 ;
   RECT 0.00 574.56 179.36 576.27 ;
   RECT 0.00 576.27 179.36 577.98 ;
   RECT 0.00 577.98 179.36 579.69 ;
   RECT 0.00 579.69 179.36 581.40 ;
   RECT 0.00 581.40 179.36 583.11 ;
   RECT 0.00 583.11 179.36 584.82 ;
   RECT 0.00 584.82 179.36 586.53 ;
   RECT 0.00 586.53 179.36 588.24 ;
   RECT 0.00 588.24 179.36 589.95 ;
   RECT 0.00 589.95 179.36 591.66 ;
   RECT 0.00 591.66 179.36 593.37 ;
   RECT 0.00 593.37 179.36 595.08 ;
   RECT 0.00 595.08 179.36 596.79 ;
   RECT 0.00 596.79 179.36 598.50 ;
   RECT 0.00 598.50 179.36 600.21 ;
   RECT 0.00 600.21 179.36 601.92 ;
   RECT 0.00 601.92 179.36 603.63 ;
   RECT 0.00 603.63 179.36 605.34 ;
   RECT 0.00 605.34 179.36 607.05 ;
   RECT 0.00 607.05 179.36 608.76 ;
   RECT 0.00 608.76 179.36 610.47 ;
   RECT 0.00 610.47 179.36 612.18 ;
   RECT 0.00 612.18 179.36 613.89 ;
   RECT 0.00 613.89 179.36 615.60 ;
   RECT 0.00 615.60 179.36 617.31 ;
   RECT 0.00 617.31 179.36 619.02 ;
   RECT 0.00 619.02 179.36 620.73 ;
   RECT 0.00 620.73 179.36 622.44 ;
   RECT 0.00 622.44 179.36 624.15 ;
   RECT 0.00 624.15 179.36 625.86 ;
   RECT 0.00 625.86 179.36 627.57 ;
   RECT 0.00 627.57 179.36 629.28 ;
   RECT 0.00 629.28 179.36 630.99 ;
   RECT 0.00 630.99 179.36 632.70 ;
   RECT 0.00 632.70 179.36 634.41 ;
   RECT 0.00 634.41 179.36 636.12 ;
   RECT 0.00 636.12 179.36 637.83 ;
   RECT 0.00 637.83 179.36 639.54 ;
   RECT 0.00 639.54 179.36 641.25 ;
   RECT 0.00 641.25 179.36 642.96 ;
   RECT 0.00 642.96 179.36 644.67 ;
   RECT 0.00 644.67 179.36 646.38 ;
   RECT 0.00 646.38 179.36 648.09 ;
   RECT 0.00 648.09 179.36 649.80 ;
   RECT 0.00 649.80 179.36 651.51 ;
   RECT 0.00 651.51 179.36 653.22 ;
   RECT 0.00 653.22 179.36 654.93 ;
   RECT 0.00 654.93 179.36 656.64 ;
   RECT 0.00 656.64 179.36 658.35 ;
   RECT 0.00 658.35 179.36 660.06 ;
   RECT 0.00 660.06 179.36 661.77 ;
   RECT 0.00 661.77 179.36 663.48 ;
   RECT 0.00 663.48 179.36 665.19 ;
   RECT 0.00 665.19 179.36 666.90 ;
   RECT 0.00 666.90 179.36 668.61 ;
   RECT 0.00 668.61 179.36 670.32 ;
   RECT 0.00 670.32 179.36 672.03 ;
   RECT 0.00 672.03 179.36 673.74 ;
   RECT 0.00 673.74 179.36 675.45 ;
   RECT 0.00 675.45 179.36 677.16 ;
   RECT 0.00 677.16 179.36 678.87 ;
   RECT 0.00 678.87 179.36 680.58 ;
   RECT 0.00 680.58 179.36 682.29 ;
   RECT 0.00 682.29 179.36 684.00 ;
   RECT 0.00 684.00 179.36 685.71 ;
   RECT 0.00 685.71 179.36 687.42 ;
   RECT 0.00 687.42 179.36 689.13 ;
   RECT 0.00 689.13 179.36 690.84 ;
   RECT 0.00 690.84 179.36 692.55 ;
   RECT 0.00 692.55 179.36 694.26 ;
   RECT 0.00 694.26 179.36 695.97 ;
   RECT 0.00 695.97 179.36 697.68 ;
   RECT 0.00 697.68 179.36 699.39 ;
   RECT 0.00 699.39 179.36 701.10 ;
   RECT 0.00 701.10 179.36 702.81 ;
   RECT 0.00 702.81 179.36 704.52 ;
   RECT 0.00 704.52 179.36 706.23 ;
   RECT 0.00 706.23 179.36 707.94 ;
   RECT 0.00 707.94 179.36 709.65 ;
   RECT 0.00 709.65 179.36 711.36 ;
   RECT 0.00 711.36 179.36 713.07 ;
   RECT 0.00 713.07 179.36 714.78 ;
   RECT 0.00 714.78 179.36 716.49 ;
   RECT 0.00 716.49 179.36 718.20 ;
   RECT 0.00 718.20 179.36 719.91 ;
   RECT 0.00 719.91 179.36 721.62 ;
   RECT 0.00 721.62 179.36 723.33 ;
   RECT 0.00 723.33 179.36 725.04 ;
   RECT 0.00 725.04 179.36 726.75 ;
   RECT 0.00 726.75 179.36 728.46 ;
   RECT 0.00 728.46 179.36 730.17 ;
   RECT 0.00 730.17 179.36 731.88 ;
   RECT 0.00 731.88 179.36 733.59 ;
   RECT 0.00 733.59 179.36 735.30 ;
   RECT 0.00 735.30 179.36 737.01 ;
   RECT 0.00 737.01 179.36 738.72 ;
   RECT 0.00 738.72 179.36 740.43 ;
   RECT 0.00 740.43 179.36 742.14 ;
   RECT 0.00 742.14 179.36 743.85 ;
   RECT 0.00 743.85 179.36 745.56 ;
   RECT 0.00 745.56 179.36 747.27 ;
   RECT 0.00 747.27 179.36 748.98 ;
   RECT 0.00 748.98 179.36 750.69 ;
   RECT 0.00 750.69 179.36 752.40 ;
   RECT 0.00 752.40 179.36 754.11 ;
   RECT 0.00 754.11 179.36 755.82 ;
   RECT 0.00 755.82 179.36 757.53 ;
   RECT 0.00 757.53 179.36 759.24 ;
   RECT 0.00 759.24 179.36 760.95 ;
   RECT 0.00 760.95 179.36 762.66 ;
   RECT 0.00 762.66 179.36 764.37 ;
   RECT 0.00 764.37 179.36 766.08 ;
   RECT 0.00 766.08 179.36 767.79 ;
   RECT 0.00 767.79 179.36 769.50 ;
   RECT 0.00 769.50 179.36 771.21 ;
   RECT 0.00 771.21 179.36 772.92 ;
   RECT 0.00 772.92 179.36 774.63 ;
   RECT 0.00 774.63 179.36 776.34 ;
   RECT 0.00 776.34 179.36 778.05 ;
   RECT 0.00 778.05 179.36 779.76 ;
   RECT 0.00 779.76 179.36 781.47 ;
   RECT 0.00 781.47 179.36 783.18 ;
   RECT 0.00 783.18 179.36 784.89 ;
   RECT 0.00 784.89 179.36 786.60 ;
   RECT 0.00 786.60 179.36 788.31 ;
   RECT 0.00 788.31 179.36 790.02 ;
   RECT 0.00 790.02 179.36 791.73 ;
   RECT 0.00 791.73 179.36 793.44 ;
   RECT 0.00 793.44 179.36 795.15 ;
   RECT 0.00 795.15 179.36 796.86 ;
   RECT 0.00 796.86 179.36 798.57 ;
   RECT 0.00 798.57 179.36 800.28 ;
   RECT 0.00 800.28 179.36 801.99 ;
   RECT 0.00 801.99 179.36 803.70 ;
   RECT 0.00 803.70 179.36 805.41 ;
   RECT 0.00 805.41 179.36 807.12 ;
   RECT 0.00 807.12 179.36 808.83 ;
   RECT 0.00 808.83 179.36 810.54 ;
   RECT 0.00 810.54 179.36 812.25 ;
   RECT 0.00 812.25 179.36 813.96 ;
   RECT 0.00 813.96 179.36 815.67 ;
   RECT 0.00 815.67 179.36 817.38 ;
   RECT 0.00 817.38 179.36 819.09 ;
   RECT 0.00 819.09 179.36 820.80 ;
   RECT 0.00 820.80 179.36 822.51 ;
   RECT 0.00 822.51 179.36 824.22 ;
   RECT 0.00 824.22 179.36 825.93 ;
   RECT 0.00 825.93 179.36 827.64 ;
   RECT 0.00 827.64 179.36 829.35 ;
   RECT 0.00 829.35 179.36 831.06 ;
   RECT 0.00 831.06 179.36 832.77 ;
   RECT 0.00 832.77 179.36 834.48 ;
   RECT 0.00 834.48 179.36 836.19 ;
   RECT 0.00 836.19 179.36 837.90 ;
   RECT 0.00 837.90 179.36 839.61 ;
   RECT 0.00 839.61 179.36 841.32 ;
 END
END block_533x4428_789f

MACRO block_416x450_106
 CLASS BLOCK ;
 FOREIGN block_416x450_106 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 158.08 BY 85.5 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 64.315 154.945 64.885 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 20.615 154.945 21.185 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 4.655 3.325 5.225 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 8.075 3.325 8.645 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 9.215 3.325 9.785 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 12.635 3.325 13.205 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 24.415 3.325 24.985 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 25.555 3.325 26.125 ;
  END
 END o7
 PIN o8
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 26.315 3.325 26.885 ;
  END
 END o8
 PIN o9
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 27.455 3.325 28.025 ;
  END
 END o9
 PIN o10
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 28.975 3.325 29.545 ;
  END
 END o10
 PIN o11
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 22.895 3.325 23.465 ;
  END
 END o11
 PIN o12
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 32.015 3.325 32.585 ;
  END
 END o12
 PIN o13
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 33.535 3.325 34.105 ;
  END
 END o13
 PIN o14
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 34.295 3.325 34.865 ;
  END
 END o14
 PIN o15
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 35.055 3.325 35.625 ;
  END
 END o15
 PIN o16
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 35.815 3.325 36.385 ;
  END
 END o16
 PIN o17
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 30.875 3.325 31.445 ;
  END
 END o17
 PIN o18
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 38.855 3.325 39.425 ;
  END
 END o18
 PIN o19
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 39.615 3.325 40.185 ;
  END
 END o19
 PIN o20
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 40.375 3.325 40.945 ;
  END
 END o20
 PIN o21
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 41.135 3.325 41.705 ;
  END
 END o21
 PIN o22
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 42.655 3.325 43.225 ;
  END
 END o22
 PIN o23
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 38.095 3.325 38.665 ;
  END
 END o23
 PIN o24
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 44.935 3.325 45.505 ;
  END
 END o24
 PIN o25
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 45.695 3.325 46.265 ;
  END
 END o25
 PIN o26
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 47.215 3.325 47.785 ;
  END
 END o26
 PIN o27
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 47.975 3.325 48.545 ;
  END
 END o27
 PIN o28
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 48.735 3.325 49.305 ;
  END
 END o28
 PIN o29
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 44.175 3.325 44.745 ;
  END
 END o29
 PIN o30
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 51.775 3.325 52.345 ;
  END
 END o30
 PIN o31
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 52.535 3.325 53.105 ;
  END
 END o31
 PIN o32
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 53.295 3.325 53.865 ;
  END
 END o32
 PIN o33
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 54.055 3.325 54.625 ;
  END
 END o33
 PIN o34
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 54.815 3.325 55.385 ;
  END
 END o34
 PIN o35
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 50.255 3.325 50.825 ;
  END
 END o35
 PIN o36
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 57.855 3.325 58.425 ;
  END
 END o36
 PIN o37
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 58.615 3.325 59.185 ;
  END
 END o37
 PIN o38
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 59.375 3.325 59.945 ;
  END
 END o38
 PIN o39
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 60.895 3.325 61.465 ;
  END
 END o39
 PIN o40
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 61.655 3.325 62.225 ;
  END
 END o40
 PIN o41
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 57.095 3.325 57.665 ;
  END
 END o41
 PIN o42
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 63.935 3.325 64.505 ;
  END
 END o42
 PIN o43
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 65.455 3.325 66.025 ;
  END
 END o43
 PIN o44
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 66.215 3.325 66.785 ;
  END
 END o44
 PIN o45
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 66.975 3.325 67.545 ;
  END
 END o45
 PIN o46
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 67.735 3.325 68.305 ;
  END
 END o46
 PIN o47
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 63.175 3.325 63.745 ;
  END
 END o47
 PIN o48
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 70.775 3.325 71.345 ;
  END
 END o48
 PIN o49
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 71.535 3.325 72.105 ;
  END
 END o49
 PIN o50
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 72.295 3.325 72.865 ;
  END
 END o50
 PIN o51
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 72.675 4.085 73.245 ;
  END
 END o51
 PIN o52
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 73.055 3.325 73.625 ;
  END
 END o52
 PIN o53
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 70.015 3.325 70.585 ;
  END
 END o53
 PIN o54
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 24.415 154.945 24.985 ;
  END
 END o54
 PIN o55
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 25.175 154.945 25.745 ;
  END
 END o55
 PIN o56
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 25.935 154.945 26.505 ;
  END
 END o56
 PIN o57
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 26.695 154.945 27.265 ;
  END
 END o57
 PIN o58
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 22.895 154.945 23.465 ;
  END
 END o58
 PIN o59
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 29.735 154.945 30.305 ;
  END
 END o59
 PIN o60
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 30.495 154.945 31.065 ;
  END
 END o60
 PIN o61
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 31.255 154.945 31.825 ;
  END
 END o61
 PIN o62
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 32.015 154.945 32.585 ;
  END
 END o62
 PIN o63
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 28.975 154.945 29.545 ;
  END
 END o63
 PIN o64
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 22.135 154.945 22.705 ;
  END
 END o64
 PIN o65
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 74.955 3.325 75.525 ;
  END
 END o65
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 51.775 154.945 52.345 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 66.975 154.945 67.545 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 49.495 154.945 50.065 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 50.255 154.945 50.825 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 54.055 154.945 54.625 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 53.295 154.945 53.865 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 47.215 154.945 47.785 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 47.975 154.945 48.545 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 3.515 3.325 4.085 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 19.855 154.945 20.425 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 18.335 154.945 18.905 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 17.575 154.945 18.145 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 48.735 154.945 49.305 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 45.695 154.945 46.265 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 44.935 154.945 45.505 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 74.575 4.085 75.145 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 21.375 154.945 21.945 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 57.095 154.945 57.665 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 57.855 154.945 58.425 ;
  END
 END i18
 PIN i19
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 58.615 154.945 59.185 ;
  END
 END i19
 PIN i20
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 59.375 154.945 59.945 ;
  END
 END i20
 PIN i21
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 60.895 154.945 61.465 ;
  END
 END i21
 PIN i22
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 61.655 154.945 62.225 ;
  END
 END i22
 PIN i23
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 62.415 154.945 62.985 ;
  END
 END i23
 PIN i24
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 63.175 154.945 63.745 ;
  END
 END i24
 PIN i25
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 3.135 154.945 3.705 ;
  END
 END i25
 PIN i26
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 3.895 154.945 4.465 ;
  END
 END i26
 PIN i27
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 4.655 154.945 5.225 ;
  END
 END i27
 PIN i28
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 6.175 154.945 6.745 ;
  END
 END i28
 PIN i29
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 6.935 154.945 7.505 ;
  END
 END i29
 PIN i30
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 7.695 154.945 8.265 ;
  END
 END i30
 PIN i31
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 8.455 154.945 9.025 ;
  END
 END i31
 PIN i32
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 9.215 154.945 9.785 ;
  END
 END i32
 PIN i33
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 10.735 154.945 11.305 ;
  END
 END i33
 PIN i34
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 11.495 154.945 12.065 ;
  END
 END i34
 PIN i35
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 12.255 154.945 12.825 ;
  END
 END i35
 PIN i36
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 13.015 154.945 13.585 ;
  END
 END i36
 PIN i37
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 13.775 154.945 14.345 ;
  END
 END i37
 PIN i38
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 15.295 154.945 15.865 ;
  END
 END i38
 PIN i39
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 16.055 154.945 16.625 ;
  END
 END i39
 OBS
  LAYER metal1 ;
   RECT 0 0 158.08 85.5 ;
  LAYER via1 ;
   RECT 0 0 158.08 85.5 ;
  LAYER metal2 ;
   RECT 0 0 158.08 85.5 ;
  LAYER via2 ;
   RECT 0 0 158.08 85.5 ;
  LAYER metal3 ;
   RECT 0 0 158.08 85.5 ;
  LAYER via3 ;
   RECT 0 0 158.08 85.5 ;
  LAYER metal4 ;
   RECT 0 0 158.08 85.5 ;
 END
END block_416x450_106

MACRO block_416x441_106
 CLASS BLOCK ;
 FOREIGN block_416x441_106 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 158.08 BY 83.79 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 64.315 154.945 64.885 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 20.615 154.945 21.185 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 4.655 3.325 5.225 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 8.075 3.325 8.645 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 9.215 3.325 9.785 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 12.635 3.325 13.205 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 24.415 3.325 24.985 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 25.555 3.325 26.125 ;
  END
 END o7
 PIN o8
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 26.315 3.325 26.885 ;
  END
 END o8
 PIN o9
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 27.455 3.325 28.025 ;
  END
 END o9
 PIN o10
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 28.975 3.325 29.545 ;
  END
 END o10
 PIN o11
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 22.895 3.325 23.465 ;
  END
 END o11
 PIN o12
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 32.015 3.325 32.585 ;
  END
 END o12
 PIN o13
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 33.535 3.325 34.105 ;
  END
 END o13
 PIN o14
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 34.295 3.325 34.865 ;
  END
 END o14
 PIN o15
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 35.055 3.325 35.625 ;
  END
 END o15
 PIN o16
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 35.815 3.325 36.385 ;
  END
 END o16
 PIN o17
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 30.875 3.325 31.445 ;
  END
 END o17
 PIN o18
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 38.855 3.325 39.425 ;
  END
 END o18
 PIN o19
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 39.615 3.325 40.185 ;
  END
 END o19
 PIN o20
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 40.375 3.325 40.945 ;
  END
 END o20
 PIN o21
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 41.135 3.325 41.705 ;
  END
 END o21
 PIN o22
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 42.655 3.325 43.225 ;
  END
 END o22
 PIN o23
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 38.095 3.325 38.665 ;
  END
 END o23
 PIN o24
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 44.935 3.325 45.505 ;
  END
 END o24
 PIN o25
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 45.695 3.325 46.265 ;
  END
 END o25
 PIN o26
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 47.215 3.325 47.785 ;
  END
 END o26
 PIN o27
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 47.975 3.325 48.545 ;
  END
 END o27
 PIN o28
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 48.735 3.325 49.305 ;
  END
 END o28
 PIN o29
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 44.175 3.325 44.745 ;
  END
 END o29
 PIN o30
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 51.775 3.325 52.345 ;
  END
 END o30
 PIN o31
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 52.535 3.325 53.105 ;
  END
 END o31
 PIN o32
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 53.295 3.325 53.865 ;
  END
 END o32
 PIN o33
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 54.055 3.325 54.625 ;
  END
 END o33
 PIN o34
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 54.815 3.325 55.385 ;
  END
 END o34
 PIN o35
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 50.255 3.325 50.825 ;
  END
 END o35
 PIN o36
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 57.855 3.325 58.425 ;
  END
 END o36
 PIN o37
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 58.615 3.325 59.185 ;
  END
 END o37
 PIN o38
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 59.375 3.325 59.945 ;
  END
 END o38
 PIN o39
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 60.895 3.325 61.465 ;
  END
 END o39
 PIN o40
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 61.655 3.325 62.225 ;
  END
 END o40
 PIN o41
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 57.095 3.325 57.665 ;
  END
 END o41
 PIN o42
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 63.935 3.325 64.505 ;
  END
 END o42
 PIN o43
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 65.455 3.325 66.025 ;
  END
 END o43
 PIN o44
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 66.215 3.325 66.785 ;
  END
 END o44
 PIN o45
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 66.975 3.325 67.545 ;
  END
 END o45
 PIN o46
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 67.735 3.325 68.305 ;
  END
 END o46
 PIN o47
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 63.175 3.325 63.745 ;
  END
 END o47
 PIN o48
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 70.775 3.325 71.345 ;
  END
 END o48
 PIN o49
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 71.535 3.325 72.105 ;
  END
 END o49
 PIN o50
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 72.295 3.325 72.865 ;
  END
 END o50
 PIN o51
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 72.675 4.085 73.245 ;
  END
 END o51
 PIN o52
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 73.055 3.325 73.625 ;
  END
 END o52
 PIN o53
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 70.015 3.325 70.585 ;
  END
 END o53
 PIN o54
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 24.415 154.945 24.985 ;
  END
 END o54
 PIN o55
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 25.175 154.945 25.745 ;
  END
 END o55
 PIN o56
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 25.935 154.945 26.505 ;
  END
 END o56
 PIN o57
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 26.695 154.945 27.265 ;
  END
 END o57
 PIN o58
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 22.895 154.945 23.465 ;
  END
 END o58
 PIN o59
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 29.735 154.945 30.305 ;
  END
 END o59
 PIN o60
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 30.495 154.945 31.065 ;
  END
 END o60
 PIN o61
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 31.255 154.945 31.825 ;
  END
 END o61
 PIN o62
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 32.015 154.945 32.585 ;
  END
 END o62
 PIN o63
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 28.975 154.945 29.545 ;
  END
 END o63
 PIN o64
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 22.135 154.945 22.705 ;
  END
 END o64
 PIN o65
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 74.955 3.325 75.525 ;
  END
 END o65
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 51.775 154.945 52.345 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 66.975 154.945 67.545 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 49.495 154.945 50.065 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 50.255 154.945 50.825 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 54.055 154.945 54.625 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 53.295 154.945 53.865 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 47.215 154.945 47.785 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 47.975 154.945 48.545 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 2.755 3.515 3.325 4.085 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 19.855 154.945 20.425 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 18.335 154.945 18.905 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 17.575 154.945 18.145 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 48.735 154.945 49.305 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 45.695 154.945 46.265 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 44.935 154.945 45.505 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 74.575 4.085 75.145 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 21.375 154.945 21.945 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 57.095 154.945 57.665 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 57.855 154.945 58.425 ;
  END
 END i18
 PIN i19
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 58.615 154.945 59.185 ;
  END
 END i19
 PIN i20
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 59.375 154.945 59.945 ;
  END
 END i20
 PIN i21
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 60.895 154.945 61.465 ;
  END
 END i21
 PIN i22
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 61.655 154.945 62.225 ;
  END
 END i22
 PIN i23
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 62.415 154.945 62.985 ;
  END
 END i23
 PIN i24
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 63.175 154.945 63.745 ;
  END
 END i24
 PIN i25
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 3.135 154.945 3.705 ;
  END
 END i25
 PIN i26
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 3.895 154.945 4.465 ;
  END
 END i26
 PIN i27
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 4.655 154.945 5.225 ;
  END
 END i27
 PIN i28
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 6.175 154.945 6.745 ;
  END
 END i28
 PIN i29
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 6.935 154.945 7.505 ;
  END
 END i29
 PIN i30
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 7.695 154.945 8.265 ;
  END
 END i30
 PIN i31
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 8.455 154.945 9.025 ;
  END
 END i31
 PIN i32
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 9.215 154.945 9.785 ;
  END
 END i32
 PIN i33
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 10.735 154.945 11.305 ;
  END
 END i33
 PIN i34
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 11.495 154.945 12.065 ;
  END
 END i34
 PIN i35
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 12.255 154.945 12.825 ;
  END
 END i35
 PIN i36
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 13.015 154.945 13.585 ;
  END
 END i36
 PIN i37
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 13.775 154.945 14.345 ;
  END
 END i37
 PIN i38
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 15.295 154.945 15.865 ;
  END
 END i38
 PIN i39
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 154.375 16.055 154.945 16.625 ;
  END
 END i39
 OBS
  LAYER metal1 ;
   RECT 0 0 158.08 83.79 ;
  LAYER via1 ;
   RECT 0 0 158.08 83.79 ;
  LAYER metal2 ;
   RECT 0 0 158.08 83.79 ;
  LAYER via2 ;
   RECT 0 0 158.08 83.79 ;
  LAYER metal3 ;
   RECT 0 0 158.08 83.79 ;
  LAYER via3 ;
   RECT 0 0 158.08 83.79 ;
  LAYER metal4 ;
   RECT 0 0 158.08 83.79 ;
 END
END block_416x441_106

MACRO block_315x2106_146
 CLASS BLOCK ;
 FOREIGN block_315x2106_146 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 119.7 BY 400.14 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 396.055 9.785 396.625 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 338.675 9.785 339.245 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 332.975 9.785 333.545 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 327.085 9.785 327.655 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 321.385 9.785 321.955 ;
  END
 END o4
 PIN o5
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 315.685 9.785 316.255 ;
  END
 END o5
 PIN o6
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 309.985 9.785 310.555 ;
  END
 END o6
 PIN o7
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 304.095 9.785 304.665 ;
  END
 END o7
 PIN o8
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 298.395 9.785 298.965 ;
  END
 END o8
 PIN o9
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 292.695 9.785 293.265 ;
  END
 END o9
 PIN o10
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 286.995 9.785 287.565 ;
  END
 END o10
 PIN o11
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 390.355 9.785 390.925 ;
  END
 END o11
 PIN o12
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 281.105 9.785 281.675 ;
  END
 END o12
 PIN o13
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 275.405 9.785 275.975 ;
  END
 END o13
 PIN o14
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 269.705 9.785 270.275 ;
  END
 END o14
 PIN o15
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 264.005 9.785 264.575 ;
  END
 END o15
 PIN o16
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 258.115 9.785 258.685 ;
  END
 END o16
 PIN o17
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 252.415 9.785 252.985 ;
  END
 END o17
 PIN o18
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 246.715 9.785 247.285 ;
  END
 END o18
 PIN o19
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 241.015 9.785 241.585 ;
  END
 END o19
 PIN o20
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 235.125 9.785 235.695 ;
  END
 END o20
 PIN o21
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 229.425 9.785 229.995 ;
  END
 END o21
 PIN o22
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 384.655 9.785 385.225 ;
  END
 END o22
 PIN o23
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 223.725 9.785 224.295 ;
  END
 END o23
 PIN o24
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 218.025 9.785 218.595 ;
  END
 END o24
 PIN o25
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 186.485 9.785 187.055 ;
  END
 END o25
 PIN o26
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 180.595 9.785 181.165 ;
  END
 END o26
 PIN o27
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 174.895 9.785 175.465 ;
  END
 END o27
 PIN o28
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 169.195 9.785 169.765 ;
  END
 END o28
 PIN o29
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 163.495 9.785 164.065 ;
  END
 END o29
 PIN o30
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 157.605 9.785 158.175 ;
  END
 END o30
 PIN o31
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 151.905 9.785 152.475 ;
  END
 END o31
 PIN o32
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 146.205 9.785 146.775 ;
  END
 END o32
 PIN o33
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 378.955 9.785 379.525 ;
  END
 END o33
 PIN o34
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 140.505 9.785 141.075 ;
  END
 END o34
 PIN o35
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 134.615 9.785 135.185 ;
  END
 END o35
 PIN o36
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 128.915 9.785 129.485 ;
  END
 END o36
 PIN o37
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 123.215 9.785 123.785 ;
  END
 END o37
 PIN o38
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 117.515 9.785 118.085 ;
  END
 END o38
 PIN o39
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 111.625 9.785 112.195 ;
  END
 END o39
 PIN o40
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 105.925 9.785 106.495 ;
  END
 END o40
 PIN o41
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 100.225 9.785 100.795 ;
  END
 END o41
 PIN o42
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 94.525 9.785 95.095 ;
  END
 END o42
 PIN o43
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 88.635 9.785 89.205 ;
  END
 END o43
 PIN o44
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 373.065 9.785 373.635 ;
  END
 END o44
 PIN o45
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 82.935 9.785 83.505 ;
  END
 END o45
 PIN o46
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 77.235 9.785 77.805 ;
  END
 END o46
 PIN o47
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 71.535 9.785 72.105 ;
  END
 END o47
 PIN o48
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 65.645 9.785 66.215 ;
  END
 END o48
 PIN o49
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 59.945 9.785 60.515 ;
  END
 END o49
 PIN o50
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 54.245 9.785 54.815 ;
  END
 END o50
 PIN o51
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 48.545 9.785 49.115 ;
  END
 END o51
 PIN o52
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 42.655 9.785 43.225 ;
  END
 END o52
 PIN o53
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 36.955 9.785 37.525 ;
  END
 END o53
 PIN o54
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 31.255 9.785 31.825 ;
  END
 END o54
 PIN o55
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 367.365 9.785 367.935 ;
  END
 END o55
 PIN o56
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 25.555 9.785 26.125 ;
  END
 END o56
 PIN o57
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 19.665 9.785 20.235 ;
  END
 END o57
 PIN o58
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 13.965 9.785 14.535 ;
  END
 END o58
 PIN o59
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 8.265 9.785 8.835 ;
  END
 END o59
 PIN o60
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 2.565 9.785 3.135 ;
  END
 END o60
 PIN o61
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 361.665 9.785 362.235 ;
  END
 END o61
 PIN o62
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 355.965 9.785 356.535 ;
  END
 END o62
 PIN o63
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 350.075 9.785 350.645 ;
  END
 END o63
 PIN o64
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 344.375 9.785 344.945 ;
  END
 END o64
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 203.585 118.465 204.155 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 195.415 118.465 195.985 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 194.085 118.465 194.655 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 111.815 194.275 112.385 194.845 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 196.935 118.465 197.505 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.135 197.505 117.705 198.075 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 195.035 9.785 195.605 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 210.995 118.465 211.565 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 200.925 118.465 201.495 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 202.255 118.465 202.825 ;
  END
 END i9
 PIN i10
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 202.065 9.785 202.635 ;
  END
 END i10
 PIN i11
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 8.455 208.715 9.025 209.285 ;
  END
 END i11
 PIN i12
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 9.215 205.675 9.785 206.245 ;
  END
 END i12
 PIN i13
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.135 203.965 117.705 204.535 ;
  END
 END i13
 PIN i14
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 205.865 118.465 206.435 ;
  END
 END i14
 PIN i15
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.135 206.245 117.705 206.815 ;
  END
 END i15
 PIN i16
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 395.675 118.465 396.245 ;
  END
 END i16
 PIN i17
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 338.295 118.465 338.865 ;
  END
 END i17
 PIN i18
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 332.405 118.465 332.975 ;
  END
 END i18
 PIN i19
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 326.705 118.465 327.275 ;
  END
 END i19
 PIN i20
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 321.005 118.465 321.575 ;
  END
 END i20
 PIN i21
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 315.305 118.465 315.875 ;
  END
 END i21
 PIN i22
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 309.415 118.465 309.985 ;
  END
 END i22
 PIN i23
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 303.715 118.465 304.285 ;
  END
 END i23
 PIN i24
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 298.015 118.465 298.585 ;
  END
 END i24
 PIN i25
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 292.315 118.465 292.885 ;
  END
 END i25
 PIN i26
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 286.425 118.465 286.995 ;
  END
 END i26
 PIN i27
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 389.975 118.465 390.545 ;
  END
 END i27
 PIN i28
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 280.725 118.465 281.295 ;
  END
 END i28
 PIN i29
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 275.025 118.465 275.595 ;
  END
 END i29
 PIN i30
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 269.325 118.465 269.895 ;
  END
 END i30
 PIN i31
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 263.435 118.465 264.005 ;
  END
 END i31
 PIN i32
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 257.735 118.465 258.305 ;
  END
 END i32
 PIN i33
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 252.035 118.465 252.605 ;
  END
 END i33
 PIN i34
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 246.335 118.465 246.905 ;
  END
 END i34
 PIN i35
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 240.445 118.465 241.015 ;
  END
 END i35
 PIN i36
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 234.745 118.465 235.315 ;
  END
 END i36
 PIN i37
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 229.045 118.465 229.615 ;
  END
 END i37
 PIN i38
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 384.275 118.465 384.845 ;
  END
 END i38
 PIN i39
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 223.345 118.465 223.915 ;
  END
 END i39
 PIN i40
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 217.455 118.465 218.025 ;
  END
 END i40
 PIN i41
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 186.865 118.465 187.435 ;
  END
 END i41
 PIN i42
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 181.165 118.465 181.735 ;
  END
 END i42
 PIN i43
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 175.275 118.465 175.845 ;
  END
 END i43
 PIN i44
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 169.575 118.465 170.145 ;
  END
 END i44
 PIN i45
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 163.875 118.465 164.445 ;
  END
 END i45
 PIN i46
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 158.175 118.465 158.745 ;
  END
 END i46
 PIN i47
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 152.285 118.465 152.855 ;
  END
 END i47
 PIN i48
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 146.585 118.465 147.155 ;
  END
 END i48
 PIN i49
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 378.385 118.465 378.955 ;
  END
 END i49
 PIN i50
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 140.885 118.465 141.455 ;
  END
 END i50
 PIN i51
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 135.185 118.465 135.755 ;
  END
 END i51
 PIN i52
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 129.295 118.465 129.865 ;
  END
 END i52
 PIN i53
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 123.595 118.465 124.165 ;
  END
 END i53
 PIN i54
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 117.895 118.465 118.465 ;
  END
 END i54
 PIN i55
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 112.195 118.465 112.765 ;
  END
 END i55
 PIN i56
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 106.305 118.465 106.875 ;
  END
 END i56
 PIN i57
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 100.605 118.465 101.175 ;
  END
 END i57
 PIN i58
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 94.905 118.465 95.475 ;
  END
 END i58
 PIN i59
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 89.205 118.465 89.775 ;
  END
 END i59
 PIN i60
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 372.685 118.465 373.255 ;
  END
 END i60
 PIN i61
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 83.315 118.465 83.885 ;
  END
 END i61
 PIN i62
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 77.615 118.465 78.185 ;
  END
 END i62
 PIN i63
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 71.915 118.465 72.485 ;
  END
 END i63
 PIN i64
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 66.215 118.465 66.785 ;
  END
 END i64
 PIN i65
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 60.325 118.465 60.895 ;
  END
 END i65
 PIN i66
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 54.625 118.465 55.195 ;
  END
 END i66
 PIN i67
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 48.925 118.465 49.495 ;
  END
 END i67
 PIN i68
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 43.225 118.465 43.795 ;
  END
 END i68
 PIN i69
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 37.335 118.465 37.905 ;
  END
 END i69
 PIN i70
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 31.635 118.465 32.205 ;
  END
 END i70
 PIN i71
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 366.985 118.465 367.555 ;
  END
 END i71
 PIN i72
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 25.935 118.465 26.505 ;
  END
 END i72
 PIN i73
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 20.235 118.465 20.805 ;
  END
 END i73
 PIN i74
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 14.345 118.465 14.915 ;
  END
 END i74
 PIN i75
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 8.645 118.465 9.215 ;
  END
 END i75
 PIN i76
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 2.945 118.465 3.515 ;
  END
 END i76
 PIN i77
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 361.285 118.465 361.855 ;
  END
 END i77
 PIN i78
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 355.395 118.465 355.965 ;
  END
 END i78
 PIN i79
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 349.695 118.465 350.265 ;
  END
 END i79
 PIN i80
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 117.895 343.995 118.465 344.565 ;
  END
 END i80
 OBS
  LAYER metal1 ;
   RECT 0 0 119.7 400.14 ;
  LAYER via1 ;
   RECT 0 0 119.7 400.14 ;
  LAYER metal2 ;
   RECT 0 0 119.7 400.14 ;
  LAYER via2 ;
   RECT 0 0 119.7 400.14 ;
  LAYER metal3 ;
   RECT 0 0 119.7 400.14 ;
  LAYER via3 ;
   RECT 0 0 119.7 400.14 ;
  LAYER metal4 ;
   RECT 0 0 119.7 400.14 ;
 END
END block_315x2106_146

MACRO block_73x72_14
 CLASS BLOCK ;
 FOREIGN block_73x72_14 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 27.74 BY 13.68 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 6.175 6.745 6.745 7.315 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 22.515 8.265 23.085 8.835 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 22.515 4.465 23.085 5.035 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 21.755 5.035 22.325 5.605 ;
  END
 END o3
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 4.275 4.085 4.845 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 19.475 11.305 20.045 11.875 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 4.275 4.845 4.845 5.415 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 5.035 4.465 5.605 5.035 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 1.425 4.085 1.995 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 2.375 4.085 2.945 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 4.275 4.085 4.845 4.655 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 8.835 4.085 9.405 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 4.275 2.565 4.845 3.135 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 6.555 4.085 7.125 ;
  END
 END i9
 OBS
  LAYER metal1 ;
   RECT 0 0 27.74 13.68 ;
  LAYER via1 ;
   RECT 0 0 27.74 13.68 ;
  LAYER metal2 ;
   RECT 0 0 27.74 13.68 ;
  LAYER via2 ;
   RECT 0 0 27.74 13.68 ;
  LAYER metal3 ;
   RECT 0 0 27.74 13.68 ;
  LAYER via3 ;
   RECT 0 0 27.74 13.68 ;
  LAYER metal4 ;
   RECT 0 0 27.74 13.68 ;
 END
END block_73x72_14

MACRO block_73x72_15
 CLASS BLOCK ;
 FOREIGN block_73x72_15 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 27.74 BY 13.68 ;
 SYMMETRY X Y ;
 PIN o0
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 1.615 4.085 2.185 ;
  END
 END o0
 PIN o1
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 6.175 6.365 6.745 6.935 ;
  END
 END o1
 PIN o2
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 22.515 4.845 23.085 5.415 ;
  END
 END o2
 PIN o3
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 22.515 8.645 23.085 9.215 ;
  END
 END o3
 PIN o4
  DIRECTION OUTPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 21.755 8.075 22.325 8.645 ;
  END
 END o4
 PIN i0
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 19.475 1.805 20.045 2.375 ;
  END
 END i0
 PIN i1
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 8.835 4.085 9.405 ;
  END
 END i1
 PIN i2
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 4.275 8.265 4.845 8.835 ;
  END
 END i2
 PIN i3
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 5.035 8.645 5.605 9.215 ;
  END
 END i3
 PIN i4
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 11.685 4.085 12.255 ;
  END
 END i4
 PIN i5
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 10.735 4.085 11.305 ;
  END
 END i5
 PIN i6
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 4.275 9.025 4.845 9.595 ;
  END
 END i6
 PIN i7
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 4.275 4.085 4.845 ;
  END
 END i7
 PIN i8
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 4.275 10.545 4.845 11.115 ;
  END
 END i8
 PIN i9
  DIRECTION INPUT ;
  USE SIGNAL ;
  PORT
   LAYER metal4 ;
   RECT 3.515 6.555 4.085 7.125 ;
  END
 END i9
 OBS
  LAYER metal1 ;
   RECT 0 0 27.74 13.68 ;
  LAYER via1 ;
   RECT 0 0 27.74 13.68 ;
  LAYER metal2 ;
   RECT 0 0 27.74 13.68 ;
  LAYER via2 ;
   RECT 0 0 27.74 13.68 ;
  LAYER metal3 ;
   RECT 0 0 27.74 13.68 ;
  LAYER via3 ;
   RECT 0 0 27.74 13.68 ;
  LAYER metal4 ;
   RECT 0 0 27.74 13.68 ;
 END
END block_73x72_15

MACRO block_7x9_0
 CLASS BLOCK ;
 FOREIGN block_7x9_0 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 2.66 BY 1.71 ;
 SYMMETRY X Y ;
 OBS
  LAYER metal1 ;
   RECT 0 0 2.66 1.71 ;
  LAYER via1 ;
   RECT 0 0 2.66 1.71 ;
  LAYER metal2 ;
   RECT 0 0 2.66 1.71 ;
  LAYER via2 ;
   RECT 0 0 2.66 1.71 ;
  LAYER metal3 ;
   RECT 0 0 2.66 1.71 ;
  LAYER via3 ;
   RECT 0 0 2.66 1.71 ;
  LAYER metal4 ;
   RECT 0 0 2.66 1.71 ;
 END
END block_7x9_0

MACRO block_100x144_0
 CLASS BLOCK ;
 FOREIGN block_100x144_0 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 38.0 BY 27.36 ;
 SYMMETRY X Y ;
 OBS
  LAYER metal1 ;
   RECT 0 0 38.0 27.36 ;
  LAYER via1 ;
   RECT 0 0 38.0 27.36 ;
  LAYER metal2 ;
   RECT 0 0 38.0 27.36 ;
  LAYER via2 ;
   RECT 0 0 38.0 27.36 ;
  LAYER metal3 ;
   RECT 0 0 38.0 27.36 ;
  LAYER via3 ;
   RECT 0 0 38.0 27.36 ;
  LAYER metal4 ;
   RECT 0 0 38.0 27.36 ;
 END
END block_100x144_0

MACRO block_26x9_0
 CLASS BLOCK ;
 FOREIGN block_26x9_0 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 9.88 BY 1.71 ;
 SYMMETRY X Y ;
 OBS
  LAYER metal1 ;
   RECT 0 0 9.88 1.71 ;
  LAYER via1 ;
   RECT 0 0 9.88 1.71 ;
  LAYER metal2 ;
   RECT 0 0 9.88 1.71 ;
  LAYER via2 ;
   RECT 0 0 9.88 1.71 ;
  LAYER metal3 ;
   RECT 0 0 9.88 1.71 ;
  LAYER via3 ;
   RECT 0 0 9.88 1.71 ;
  LAYER metal4 ;
   RECT 0 0 9.88 1.71 ;
 END
END block_26x9_0

MACRO block_43x63_0
 CLASS BLOCK ;
 FOREIGN block_43x63_0 0.000 0.000 ;
 ORIGIN 0.000 0.000 ;
   SIZE 16.34 BY 11.97 ;
 SYMMETRY X Y ;
 OBS
  LAYER metal1 ;
   RECT 0 0 16.34 11.97 ;
  LAYER via1 ;
   RECT 0 0 16.34 11.97 ;
  LAYER metal2 ;
   RECT 0 0 16.34 11.97 ;
  LAYER via2 ;
   RECT 0 0 16.34 11.97 ;
  LAYER metal3 ;
   RECT 0 0 16.34 11.97 ;
  LAYER via3 ;
   RECT 0 0 16.34 11.97 ;
  LAYER metal4 ;
   RECT 0 0 16.34 11.97 ;
 END
END block_43x63_0

END LIBRARY
